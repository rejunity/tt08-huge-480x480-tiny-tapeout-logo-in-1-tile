/*
 * Copyright (c) 2024 Tiny Tapeout LTD
 * SPDX-License-Identifier: Apache-2.0
 * Author: Renaldas Zioma
 */

`default_nettype none

parameter LOGO_SIZE = 128;  // Size of the logo in pixels
parameter DISPLAY_WIDTH = 640;  // VGA display width
parameter DISPLAY_HEIGHT = 480;  // VGA display height

`define COLOR_WHITE 3'd7

module tt_um_rejunity_vga_logo (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // VGA signals
  wire hsync;
  wire vsync;
  reg [1:0] R;
  reg [1:0] G;
  reg [1:0] B;
  wire video_active;
  wire [9:0] pix_x;
  wire [9:0] pix_y;


  // TinyVGA PMOD
  assign uo_out  = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

  // Unused outputs assigned to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in[7:1], uio_in};

  hvsync_generator vga_sync_gen (
      .clk(clk),
      .reset(~rst_n),
      .hsync(hsync),
      .vsync(vsync),
      .display_on(video_active),
      .hpos(pix_x),
      .vpos(pix_y)
  );

  reg pixel_value;

  // bitmap_rom rom1 (
  //     .x(pix_x[6:0]),
  //     .y(pix_y[6:0]),
  //     .pixel(pixel_value)
  // );

  reg [11:0] addr;
  reg [7:0] len;
  bitmap_rom_rle rom2 (
    .addr(addr),
    .len(len)
  );

  assign {R, G, B } = video_active*pixel_value*6'b11_11_00;

  // increase couner every frame (vsync happens once per frame)
  reg [11:0] counter;
  always @(posedge clk) begin
    if (~rst_n) begin
      counter <= 0;
    end else begin
      if (vsync) begin
        addr <= 0;
        counter <= 0;
        pixel_value <= 0;
      end else if (pix_x < 272 && pix_y < 267) begin
        if (counter >= len) begin
          addr <= addr + 1;
          counter <= 0;
          pixel_value <= ~pixel_value;
        end else
          counter <= counter + 1;
      end
    end
  end  

endmodule

// --------------------------------------------------------

module bitmap_rom_rle (
    input wire [11:0] addr,
    output wire [7:0] len
);

  reg [7:0] mem[1329:0];
  initial begin
    mem[12'h0000] = 8'h87;
    mem[12'h0001] = 8'h01;
    mem[12'h0002] = 8'hfd;
    mem[12'h0003] = 8'h21;
    mem[12'h0004] = 8'he7;
    mem[12'h0005] = 8'h2d;
    mem[12'h0006] = 8'hdc;
    mem[12'h0007] = 8'h38;
    mem[12'h0008] = 8'hd1;
    mem[12'h0009] = 8'h41;
    mem[12'h000a] = 8'hca;
    mem[12'h000b] = 8'h48;
    mem[12'h000c] = 8'hc2;
    mem[12'h000d] = 8'h4f;
    mem[12'h000e] = 8'hbc;
    mem[12'h000f] = 8'h55;
    mem[12'h0010] = 8'hb6;
    mem[12'h0011] = 8'h5b;
    mem[12'h0012] = 8'hb0;
    mem[12'h0013] = 8'h61;
    mem[12'h0014] = 8'hab;
    mem[12'h0015] = 8'h65;
    mem[12'h0016] = 8'ha7;
    mem[12'h0017] = 8'h69;
    mem[12'h0018] = 8'ha2;
    mem[12'h0019] = 8'h6f;
    mem[12'h001a] = 8'h9d;
    mem[12'h001b] = 8'h73;
    mem[12'h001c] = 8'h99;
    mem[12'h001d] = 8'h77;
    mem[12'h001e] = 8'h95;
    mem[12'h001f] = 8'h7b;
    mem[12'h0020] = 8'h91;
    mem[12'h0021] = 8'h7f;
    mem[12'h0022] = 8'h8e;
    mem[12'h0023] = 8'h82;
    mem[12'h0024] = 8'h8a;
    mem[12'h0025] = 8'h85;
    mem[12'h0026] = 8'h87;
    mem[12'h0027] = 8'h89;
    mem[12'h0028] = 8'h84;
    mem[12'h0029] = 8'h8c;
    mem[12'h002a] = 8'h80;
    mem[12'h002b] = 8'h8f;
    mem[12'h002c] = 8'h7d;
    mem[12'h002d] = 8'h3c;
    mem[12'h002e] = 8'h19;
    mem[12'h002f] = 8'h3c;
    mem[12'h0030] = 8'h7a;
    mem[12'h0031] = 8'h37;
    mem[12'h0032] = 8'h25;
    mem[12'h0033] = 8'h37;
    mem[12'h0034] = 8'h77;
    mem[12'h0035] = 8'h34;
    mem[12'h0036] = 8'h2f;
    mem[12'h0037] = 8'h34;
    mem[12'h0038] = 8'h74;
    mem[12'h0039] = 8'h31;
    mem[12'h003a] = 8'h38;
    mem[12'h003b] = 8'h30;
    mem[12'h003c] = 8'h72;
    mem[12'h003d] = 8'h2e;
    mem[12'h003e] = 8'h3f;
    mem[12'h003f] = 8'h2e;
    mem[12'h0040] = 8'h6f;
    mem[12'h0041] = 8'h2d;
    mem[12'h0042] = 8'h45;
    mem[12'h0043] = 8'h2d;
    mem[12'h0044] = 8'h6c;
    mem[12'h0045] = 8'h2b;
    mem[12'h0046] = 8'h4b;
    mem[12'h0047] = 8'h2b;
    mem[12'h0048] = 8'h6a;
    mem[12'h0049] = 8'h29;
    mem[12'h004a] = 8'h51;
    mem[12'h004b] = 8'h29;
    mem[12'h004c] = 8'h68;
    mem[12'h004d] = 8'h28;
    mem[12'h004e] = 8'h55;
    mem[12'h004f] = 8'h29;
    mem[12'h0050] = 8'h64;
    mem[12'h0051] = 8'h28;
    mem[12'h0052] = 8'h59;
    mem[12'h0053] = 8'h28;
    mem[12'h0054] = 8'h62;
    mem[12'h0055] = 8'h27;
    mem[12'h0056] = 8'h5e;
    mem[12'h0057] = 8'h26;
    mem[12'h0058] = 8'h60;
    mem[12'h0059] = 8'h25;
    mem[12'h005a] = 8'h63;
    mem[12'h005b] = 8'h25;
    mem[12'h005c] = 8'h5e;
    mem[12'h005d] = 8'h24;
    mem[12'h005e] = 8'h67;
    mem[12'h005f] = 8'h24;
    mem[12'h0060] = 8'h5c;
    mem[12'h0061] = 8'h24;
    mem[12'h0062] = 8'h6a;
    mem[12'h0063] = 8'h23;
    mem[12'h0064] = 8'h5a;
    mem[12'h0065] = 8'h23;
    mem[12'h0066] = 8'h6d;
    mem[12'h0067] = 8'h23;
    mem[12'h0068] = 8'h58;
    mem[12'h0069] = 8'h22;
    mem[12'h006a] = 8'h71;
    mem[12'h006b] = 8'h23;
    mem[12'h006c] = 8'h55;
    mem[12'h006d] = 8'h21;
    mem[12'h006e] = 8'h75;
    mem[12'h006f] = 8'h22;
    mem[12'h0070] = 8'h53;
    mem[12'h0071] = 8'h21;
    mem[12'h0072] = 8'h77;
    mem[12'h0073] = 8'h22;
    mem[12'h0074] = 8'h51;
    mem[12'h0075] = 8'h20;
    mem[12'h0076] = 8'h7b;
    mem[12'h0077] = 8'h21;
    mem[12'h0078] = 8'h4f;
    mem[12'h0079] = 8'h20;
    mem[12'h007a] = 8'h7d;
    mem[12'h007b] = 8'h21;
    mem[12'h007c] = 8'h4d;
    mem[12'h007d] = 8'h1f;
    mem[12'h007e] = 8'h81;
    mem[12'h007f] = 8'h1f;
    mem[12'h0080] = 8'h4c;
    mem[12'h0081] = 8'h1f;
    mem[12'h0082] = 8'h83;
    mem[12'h0083] = 8'h1f;
    mem[12'h0084] = 8'h4a;
    mem[12'h0085] = 8'h1f;
    mem[12'h0086] = 8'h85;
    mem[12'h0087] = 8'h1f;
    mem[12'h0088] = 8'h48;
    mem[12'h0089] = 8'h1e;
    mem[12'h008a] = 8'h89;
    mem[12'h008b] = 8'h1e;
    mem[12'h008c] = 8'h46;
    mem[12'h008d] = 8'h1e;
    mem[12'h008e] = 8'h8b;
    mem[12'h008f] = 8'h1e;
    mem[12'h0090] = 8'h44;
    mem[12'h0091] = 8'h1e;
    mem[12'h0092] = 8'h8d;
    mem[12'h0093] = 8'h1e;
    mem[12'h0094] = 8'h42;
    mem[12'h0095] = 8'h1e;
    mem[12'h0096] = 8'h8f;
    mem[12'h0097] = 8'h1e;
    mem[12'h0098] = 8'h40;
    mem[12'h0099] = 8'h1d;
    mem[12'h009a] = 8'h93;
    mem[12'h009b] = 8'h1d;
    mem[12'h009c] = 8'h3f;
    mem[12'h009d] = 8'h1c;
    mem[12'h009e] = 8'h95;
    mem[12'h009f] = 8'h1c;
    mem[12'h00a0] = 8'h3e;
    mem[12'h00a1] = 8'h1c;
    mem[12'h00a2] = 8'h97;
    mem[12'h00a3] = 8'h1c;
    mem[12'h00a4] = 8'h3c;
    mem[12'h00a5] = 8'h1c;
    mem[12'h00a6] = 8'h99;
    mem[12'h00a7] = 8'h1c;
    mem[12'h00a8] = 8'h3a;
    mem[12'h00a9] = 8'h1c;
    mem[12'h00aa] = 8'h9b;
    mem[12'h00ab] = 8'h1c;
    mem[12'h00ac] = 8'h39;
    mem[12'h00ad] = 8'h1b;
    mem[12'h00ae] = 8'h9d;
    mem[12'h00af] = 8'h1c;
    mem[12'h00b0] = 8'h37;
    mem[12'h00b1] = 8'h1b;
    mem[12'h00b2] = 8'h9f;
    mem[12'h00b3] = 8'h1b;
    mem[12'h00b4] = 8'h36;
    mem[12'h00b5] = 8'h86;
    mem[12'h00b6] = 8'h36;
    mem[12'h00b7] = 8'h1b;
    mem[12'h00b8] = 8'h34;
    mem[12'h00b9] = 8'h87;
    mem[12'h00ba] = 8'h37;
    mem[12'h00bb] = 8'h1b;
    mem[12'h00bc] = 8'h33;
    mem[12'h00bd] = 8'h87;
    mem[12'h00be] = 8'h38;
    mem[12'h00bf] = 8'h1a;
    mem[12'h00c0] = 8'h32;
    mem[12'h00c1] = 8'h88;
    mem[12'h00c2] = 8'h39;
    mem[12'h00c3] = 8'h1a;
    mem[12'h00c4] = 8'h30;
    mem[12'h00c5] = 8'h89;
    mem[12'h00c6] = 8'h3a;
    mem[12'h00c7] = 8'h1a;
    mem[12'h00c8] = 8'h2f;
    mem[12'h00c9] = 8'h89;
    mem[12'h00ca] = 8'h3a;
    mem[12'h00cb] = 8'h1a;
    mem[12'h00cc] = 8'h2e;
    mem[12'h00cd] = 8'h8a;
    mem[12'h00ce] = 8'h3b;
    mem[12'h00cf] = 8'h1a;
    mem[12'h00d0] = 8'h2c;
    mem[12'h00d1] = 8'h8b;
    mem[12'h00d2] = 8'h3c;
    mem[12'h00d3] = 8'h1a;
    mem[12'h00d4] = 8'h2b;
    mem[12'h00d5] = 8'h8b;
    mem[12'h00d6] = 8'h3d;
    mem[12'h00d7] = 8'h19;
    mem[12'h00d8] = 8'h2a;
    mem[12'h00d9] = 8'h8c;
    mem[12'h00da] = 8'h3e;
    mem[12'h00db] = 8'h19;
    mem[12'h00dc] = 8'h29;
    mem[12'h00dd] = 8'h8c;
    mem[12'h00de] = 8'h3e;
    mem[12'h00df] = 8'h19;
    mem[12'h00e0] = 8'h28;
    mem[12'h00e1] = 8'h8d;
    mem[12'h00e2] = 8'h3f;
    mem[12'h00e3] = 8'h19;
    mem[12'h00e4] = 8'h27;
    mem[12'h00e5] = 8'h8d;
    mem[12'h00e6] = 8'h40;
    mem[12'h00e7] = 8'h19;
    mem[12'h00e8] = 8'h25;
    mem[12'h00e9] = 8'h8e;
    mem[12'h00ea] = 8'h41;
    mem[12'h00eb] = 8'h18;
    mem[12'h00ec] = 8'h24;
    mem[12'h00ed] = 8'h8f;
    mem[12'h00ee] = 8'h41;
    mem[12'h00ef] = 8'h19;
    mem[12'h00f0] = 8'h23;
    mem[12'h00f1] = 8'h8f;
    mem[12'h00f2] = 8'h42;
    mem[12'h00f3] = 8'h18;
    mem[12'h00f4] = 8'h22;
    mem[12'h00f5] = 8'h90;
    mem[12'h00f6] = 8'h43;
    mem[12'h00f7] = 8'h18;
    mem[12'h00f8] = 8'h21;
    mem[12'h00f9] = 8'h90;
    mem[12'h00fa] = 8'h43;
    mem[12'h00fb] = 8'h18;
    mem[12'h00fc] = 8'h20;
    mem[12'h00fd] = 8'h91;
    mem[12'h00fe] = 8'h44;
    mem[12'h00ff] = 8'h18;
    mem[12'h0100] = 8'h1f;
    mem[12'h0101] = 8'h91;
    mem[12'h0102] = 8'h45;
    mem[12'h0103] = 8'h17;
    mem[12'h0104] = 8'h1e;
    mem[12'h0105] = 8'h92;
    mem[12'h0106] = 8'h45;
    mem[12'h0107] = 8'h18;
    mem[12'h0108] = 8'h1d;
    mem[12'h0109] = 8'h92;
    mem[12'h010a] = 8'h46;
    mem[12'h010b] = 8'h17;
    mem[12'h010c] = 8'h1c;
    mem[12'h010d] = 8'h93;
    mem[12'h010e] = 8'h46;
    mem[12'h010f] = 8'h18;
    mem[12'h0110] = 8'h1b;
    mem[12'h0111] = 8'h93;
    mem[12'h0112] = 8'h47;
    mem[12'h0113] = 8'h17;
    mem[12'h0114] = 8'h1b;
    mem[12'h0115] = 8'h93;
    mem[12'h0116] = 8'h48;
    mem[12'h0117] = 8'h17;
    mem[12'h0118] = 8'h19;
    mem[12'h0119] = 8'h94;
    mem[12'h011a] = 8'h48;
    mem[12'h011b] = 8'h17;
    mem[12'h011c] = 8'h19;
    mem[12'h011d] = 8'h94;
    mem[12'h011e] = 8'h49;
    mem[12'h011f] = 8'h16;
    mem[12'h0120] = 8'h18;
    mem[12'h0121] = 8'h95;
    mem[12'h0122] = 8'h49;
    mem[12'h0123] = 8'h17;
    mem[12'h0124] = 8'h17;
    mem[12'h0125] = 8'h95;
    mem[12'h0126] = 8'h4a;
    mem[12'h0127] = 8'h16;
    mem[12'h0128] = 8'h16;
    mem[12'h0129] = 8'h96;
    mem[12'h012a] = 8'h4a;
    mem[12'h012b] = 8'h17;
    mem[12'h012c] = 8'h15;
    mem[12'h012d] = 8'h96;
    mem[12'h012e] = 8'h4b;
    mem[12'h012f] = 8'h16;
    mem[12'h0130] = 8'h15;
    mem[12'h0131] = 8'h96;
    mem[12'h0132] = 8'h4b;
    mem[12'h0133] = 8'h16;
    mem[12'h0134] = 8'h14;
    mem[12'h0135] = 8'h97;
    mem[12'h0136] = 8'h4c;
    mem[12'h0137] = 8'h16;
    mem[12'h0138] = 8'h13;
    mem[12'h0139] = 8'h97;
    mem[12'h013a] = 8'h4c;
    mem[12'h013b] = 8'h16;
    mem[12'h013c] = 8'h13;
    mem[12'h013d] = 8'h97;
    mem[12'h013e] = 8'h4c;
    mem[12'h013f] = 8'h16;
    mem[12'h0140] = 8'h12;
    mem[12'h0141] = 8'h98;
    mem[12'h0142] = 8'h4d;
    mem[12'h0143] = 8'h16;
    mem[12'h0144] = 8'h11;
    mem[12'h0145] = 8'h98;
    mem[12'h0146] = 8'h4d;
    mem[12'h0147] = 8'h16;
    mem[12'h0148] = 8'h5b;
    mem[12'h0149] = 8'h27;
    mem[12'h014a] = 8'h75;
    mem[12'h014b] = 8'h16;
    mem[12'h014c] = 8'h5a;
    mem[12'h014d] = 8'h27;
    mem[12'h014e] = 8'h75;
    mem[12'h014f] = 8'h16;
    mem[12'h0150] = 8'h5a;
    mem[12'h0151] = 8'h27;
    mem[12'h0152] = 8'h75;
    mem[12'h0153] = 8'h16;
    mem[12'h0154] = 8'h5a;
    mem[12'h0155] = 8'h27;
    mem[12'h0156] = 8'h76;
    mem[12'h0157] = 8'h15;
    mem[12'h0158] = 8'h5a;
    mem[12'h0159] = 8'h27;
    mem[12'h015a] = 8'h76;
    mem[12'h015b] = 8'h16;
    mem[12'h015c] = 8'h59;
    mem[12'h015d] = 8'h27;
    mem[12'h015e] = 8'h76;
    mem[12'h015f] = 8'h16;
    mem[12'h0160] = 8'h59;
    mem[12'h0161] = 8'h27;
    mem[12'h0162] = 8'h77;
    mem[12'h0163] = 8'h15;
    mem[12'h0164] = 8'h59;
    mem[12'h0165] = 8'h27;
    mem[12'h0166] = 8'h77;
    mem[12'h0167] = 8'h16;
    mem[12'h0168] = 8'h58;
    mem[12'h0169] = 8'h27;
    mem[12'h016a] = 8'h77;
    mem[12'h016b] = 8'h16;
    mem[12'h016c] = 8'h58;
    mem[12'h016d] = 8'h27;
    mem[12'h016e] = 8'h78;
    mem[12'h016f] = 8'h15;
    mem[12'h0170] = 8'h58;
    mem[12'h0171] = 8'h27;
    mem[12'h0172] = 8'h78;
    mem[12'h0173] = 8'h15;
    mem[12'h0174] = 8'h0b;
    mem[12'h0175] = 8'h15;
    mem[12'h0176] = 8'h36;
    mem[12'h0177] = 8'h27;
    mem[12'h0178] = 8'h78;
    mem[12'h0179] = 8'h15;
    mem[12'h017a] = 8'h0a;
    mem[12'h017b] = 8'h16;
    mem[12'h017c] = 8'h36;
    mem[12'h017d] = 8'h27;
    mem[12'h017e] = 8'h79;
    mem[12'h017f] = 8'h15;
    mem[12'h0180] = 8'h09;
    mem[12'h0181] = 8'h15;
    mem[12'h0182] = 8'h37;
    mem[12'h0183] = 8'h27;
    mem[12'h0184] = 8'h79;
    mem[12'h0185] = 8'h15;
    mem[12'h0186] = 8'h09;
    mem[12'h0187] = 8'h15;
    mem[12'h0188] = 8'h37;
    mem[12'h0189] = 8'h27;
    mem[12'h018a] = 8'h79;
    mem[12'h018b] = 8'h15;
    mem[12'h018c] = 8'h09;
    mem[12'h018d] = 8'h15;
    mem[12'h018e] = 8'h37;
    mem[12'h018f] = 8'h27;
    mem[12'h0190] = 8'h79;
    mem[12'h0191] = 8'h15;
    mem[12'h0192] = 8'h09;
    mem[12'h0193] = 8'h15;
    mem[12'h0194] = 8'h37;
    mem[12'h0195] = 8'h27;
    mem[12'h0196] = 8'h7a;
    mem[12'h0197] = 8'h14;
    mem[12'h0198] = 8'h08;
    mem[12'h0199] = 8'h15;
    mem[12'h019a] = 8'h38;
    mem[12'h019b] = 8'h27;
    mem[12'h019c] = 8'h7a;
    mem[12'h019d] = 8'h15;
    mem[12'h019e] = 8'h07;
    mem[12'h019f] = 8'h15;
    mem[12'h01a0] = 8'h38;
    mem[12'h01a1] = 8'h27;
    mem[12'h01a2] = 8'h7a;
    mem[12'h01a3] = 8'h15;
    mem[12'h01a4] = 8'h07;
    mem[12'h01a5] = 8'h15;
    mem[12'h01a6] = 8'h38;
    mem[12'h01a7] = 8'h27;
    mem[12'h01a8] = 8'h7a;
    mem[12'h01a9] = 8'h15;
    mem[12'h01aa] = 8'h07;
    mem[12'h01ab] = 8'h15;
    mem[12'h01ac] = 8'h38;
    mem[12'h01ad] = 8'h27;
    mem[12'h01ae] = 8'h7a;
    mem[12'h01af] = 8'h15;
    mem[12'h01b0] = 8'h07;
    mem[12'h01b1] = 8'h15;
    mem[12'h01b2] = 8'h38;
    mem[12'h01b3] = 8'h27;
    mem[12'h01b4] = 8'h7b;
    mem[12'h01b5] = 8'h14;
    mem[12'h01b6] = 8'h07;
    mem[12'h01b7] = 8'h14;
    mem[12'h01b8] = 8'h39;
    mem[12'h01b9] = 8'h27;
    mem[12'h01ba] = 8'h7b;
    mem[12'h01bb] = 8'h14;
    mem[12'h01bc] = 8'h06;
    mem[12'h01bd] = 8'h15;
    mem[12'h01be] = 8'h39;
    mem[12'h01bf] = 8'h27;
    mem[12'h01c0] = 8'h7b;
    mem[12'h01c1] = 8'h15;
    mem[12'h01c2] = 8'h05;
    mem[12'h01c3] = 8'h15;
    mem[12'h01c4] = 8'h39;
    mem[12'h01c5] = 8'h27;
    mem[12'h01c6] = 8'h7b;
    mem[12'h01c7] = 8'h15;
    mem[12'h01c8] = 8'h05;
    mem[12'h01c9] = 8'h15;
    mem[12'h01ca] = 8'h39;
    mem[12'h01cb] = 8'h27;
    mem[12'h01cc] = 8'h7b;
    mem[12'h01cd] = 8'h15;
    mem[12'h01ce] = 8'h05;
    mem[12'h01cf] = 8'h15;
    mem[12'h01d0] = 8'h39;
    mem[12'h01d1] = 8'h27;
    mem[12'h01d2] = 8'h7b;
    mem[12'h01d3] = 8'h15;
    mem[12'h01d4] = 8'h05;
    mem[12'h01d5] = 8'h15;
    mem[12'h01d6] = 8'h39;
    mem[12'h01d7] = 8'h27;
    mem[12'h01d8] = 8'h7b;
    mem[12'h01d9] = 8'h15;
    mem[12'h01da] = 8'h05;
    mem[12'h01db] = 8'h14;
    mem[12'h01dc] = 8'h3a;
    mem[12'h01dd] = 8'h27;
    mem[12'h01de] = 8'h7c;
    mem[12'h01df] = 8'h14;
    mem[12'h01e0] = 8'h05;
    mem[12'h01e1] = 8'h14;
    mem[12'h01e2] = 8'h3a;
    mem[12'h01e3] = 8'h8c;
    mem[12'h01e4] = 8'h17;
    mem[12'h01e5] = 8'h14;
    mem[12'h01e6] = 8'h05;
    mem[12'h01e7] = 8'h14;
    mem[12'h01e8] = 8'h3a;
    mem[12'h01e9] = 8'h8c;
    mem[12'h01ea] = 8'h17;
    mem[12'h01eb] = 8'h14;
    mem[12'h01ec] = 8'h05;
    mem[12'h01ed] = 8'h14;
    mem[12'h01ee] = 8'h3a;
    mem[12'h01ef] = 8'h8c;
    mem[12'h01f0] = 8'h17;
    mem[12'h01f1] = 8'h14;
    mem[12'h01f2] = 8'h05;
    mem[12'h01f3] = 8'h14;
    mem[12'h01f4] = 8'h3a;
    mem[12'h01f5] = 8'h8c;
    mem[12'h01f6] = 8'h17;
    mem[12'h01f7] = 8'h14;
    mem[12'h01f8] = 8'h05;
    mem[12'h01f9] = 8'h14;
    mem[12'h01fa] = 8'h3a;
    mem[12'h01fb] = 8'h8c;
    mem[12'h01fc] = 8'h17;
    mem[12'h01fd] = 8'h15;
    mem[12'h01fe] = 8'h04;
    mem[12'h01ff] = 8'h14;
    mem[12'h0200] = 8'h3a;
    mem[12'h0201] = 8'h8c;
    mem[12'h0202] = 8'h17;
    mem[12'h0203] = 8'h15;
    mem[12'h0204] = 8'h04;
    mem[12'h0205] = 8'h14;
    mem[12'h0206] = 8'h3a;
    mem[12'h0207] = 8'h8c;
    mem[12'h0208] = 8'h17;
    mem[12'h0209] = 8'h15;
    mem[12'h020a] = 8'h03;
    mem[12'h020b] = 8'h15;
    mem[12'h020c] = 8'h3a;
    mem[12'h020d] = 8'h8c;
    mem[12'h020e] = 8'h17;
    mem[12'h020f] = 8'h15;
    mem[12'h0210] = 8'h03;
    mem[12'h0211] = 8'h15;
    mem[12'h0212] = 8'h3a;
    mem[12'h0213] = 8'h8c;
    mem[12'h0214] = 8'h17;
    mem[12'h0215] = 8'h15;
    mem[12'h0216] = 8'h03;
    mem[12'h0217] = 8'h15;
    mem[12'h0218] = 8'h3a;
    mem[12'h0219] = 8'h8c;
    mem[12'h021a] = 8'h17;
    mem[12'h021b] = 8'h15;
    mem[12'h021c] = 8'h03;
    mem[12'h021d] = 8'h15;
    mem[12'h021e] = 8'h3a;
    mem[12'h021f] = 8'h8c;
    mem[12'h0220] = 8'h17;
    mem[12'h0221] = 8'h15;
    mem[12'h0222] = 8'h03;
    mem[12'h0223] = 8'h15;
    mem[12'h0224] = 8'h3a;
    mem[12'h0225] = 8'h8c;
    mem[12'h0226] = 8'h17;
    mem[12'h0227] = 8'h15;
    mem[12'h0228] = 8'h03;
    mem[12'h0229] = 8'h15;
    mem[12'h022a] = 8'h3a;
    mem[12'h022b] = 8'h8c;
    mem[12'h022c] = 8'h17;
    mem[12'h022d] = 8'h15;
    mem[12'h022e] = 8'h03;
    mem[12'h022f] = 8'h15;
    mem[12'h0230] = 8'h3a;
    mem[12'h0231] = 8'h8c;
    mem[12'h0232] = 8'h17;
    mem[12'h0233] = 8'h15;
    mem[12'h0234] = 8'h03;
    mem[12'h0235] = 8'h15;
    mem[12'h0236] = 8'h3a;
    mem[12'h0237] = 8'h8c;
    mem[12'h0238] = 8'h17;
    mem[12'h0239] = 8'h15;
    mem[12'h023a] = 8'h03;
    mem[12'h023b] = 8'h15;
    mem[12'h023c] = 8'h3a;
    mem[12'h023d] = 8'h8c;
    mem[12'h023e] = 8'h17;
    mem[12'h023f] = 8'h15;
    mem[12'h0240] = 8'h03;
    mem[12'h0241] = 8'h15;
    mem[12'h0242] = 8'h3a;
    mem[12'h0243] = 8'h8c;
    mem[12'h0244] = 8'h17;
    mem[12'h0245] = 8'h15;
    mem[12'h0246] = 8'h03;
    mem[12'h0247] = 8'h15;
    mem[12'h0248] = 8'h3a;
    mem[12'h0249] = 8'h8c;
    mem[12'h024a] = 8'h17;
    mem[12'h024b] = 8'h15;
    mem[12'h024c] = 8'h04;
    mem[12'h024d] = 8'h14;
    mem[12'h024e] = 8'h3a;
    mem[12'h024f] = 8'h8c;
    mem[12'h0250] = 8'h17;
    mem[12'h0251] = 8'h15;
    mem[12'h0252] = 8'h04;
    mem[12'h0253] = 8'h14;
    mem[12'h0254] = 8'h3a;
    mem[12'h0255] = 8'h8c;
    mem[12'h0256] = 8'h17;
    mem[12'h0257] = 8'h15;
    mem[12'h0258] = 8'h04;
    mem[12'h0259] = 8'h14;
    mem[12'h025a] = 8'h3a;
    mem[12'h025b] = 8'h8c;
    mem[12'h025c] = 8'h17;
    mem[12'h025d] = 8'h14;
    mem[12'h025e] = 8'h05;
    mem[12'h025f] = 8'h14;
    mem[12'h0260] = 8'h3a;
    mem[12'h0261] = 8'h8c;
    mem[12'h0262] = 8'h17;
    mem[12'h0263] = 8'h14;
    mem[12'h0264] = 8'h05;
    mem[12'h0265] = 8'h14;
    mem[12'h0266] = 8'h3a;
    mem[12'h0267] = 8'h8c;
    mem[12'h0268] = 8'h17;
    mem[12'h0269] = 8'h14;
    mem[12'h026a] = 8'h05;
    mem[12'h026b] = 8'h14;
    mem[12'h026c] = 8'h3a;
    mem[12'h026d] = 8'h8c;
    mem[12'h026e] = 8'h17;
    mem[12'h026f] = 8'h14;
    mem[12'h0270] = 8'h05;
    mem[12'h0271] = 8'h14;
    mem[12'h0272] = 8'h3a;
    mem[12'h0273] = 8'h8c;
    mem[12'h0274] = 8'h17;
    mem[12'h0275] = 8'h14;
    mem[12'h0276] = 8'h05;
    mem[12'h0277] = 8'h15;
    mem[12'h0278] = 8'h39;
    mem[12'h0279] = 8'h8c;
    mem[12'h027a] = 8'h17;
    mem[12'h027b] = 8'h14;
    mem[12'h027c] = 8'h05;
    mem[12'h027d] = 8'h15;
    mem[12'h027e] = 8'h39;
    mem[12'h027f] = 8'h8c;
    mem[12'h0280] = 8'h16;
    mem[12'h0281] = 8'h15;
    mem[12'h0282] = 8'h05;
    mem[12'h0283] = 8'h15;
    mem[12'h0284] = 8'h39;
    mem[12'h0285] = 8'h8c;
    mem[12'h0286] = 8'h16;
    mem[12'h0287] = 8'h15;
    mem[12'h0288] = 8'h05;
    mem[12'h0289] = 8'h15;
    mem[12'h028a] = 8'h39;
    mem[12'h028b] = 8'h8c;
    mem[12'h028c] = 8'h16;
    mem[12'h028d] = 8'h15;
    mem[12'h028e] = 8'h05;
    mem[12'h028f] = 8'h15;
    mem[12'h0290] = 8'h39;
    mem[12'h0291] = 8'h8c;
    mem[12'h0292] = 8'h16;
    mem[12'h0293] = 8'h15;
    mem[12'h0294] = 8'h06;
    mem[12'h0295] = 8'h14;
    mem[12'h0296] = 8'h39;
    mem[12'h0297] = 8'h8c;
    mem[12'h0298] = 8'h16;
    mem[12'h0299] = 8'h15;
    mem[12'h029a] = 8'h06;
    mem[12'h029b] = 8'h14;
    mem[12'h029c] = 8'h39;
    mem[12'h029d] = 8'h8c;
    mem[12'h029e] = 8'h16;
    mem[12'h029f] = 8'h14;
    mem[12'h02a0] = 8'h07;
    mem[12'h02a1] = 8'h15;
    mem[12'h02a2] = 8'h38;
    mem[12'h02a3] = 8'h8c;
    mem[12'h02a4] = 8'h15;
    mem[12'h02a5] = 8'h15;
    mem[12'h02a6] = 8'h07;
    mem[12'h02a7] = 8'h15;
    mem[12'h02a8] = 8'h38;
    mem[12'h02a9] = 8'h8c;
    mem[12'h02aa] = 8'h15;
    mem[12'h02ab] = 8'h15;
    mem[12'h02ac] = 8'h07;
    mem[12'h02ad] = 8'h15;
    mem[12'h02ae] = 8'h38;
    mem[12'h02af] = 8'h8c;
    mem[12'h02b0] = 8'h15;
    mem[12'h02b1] = 8'h15;
    mem[12'h02b2] = 8'h07;
    mem[12'h02b3] = 8'h15;
    mem[12'h02b4] = 8'h38;
    mem[12'h02b5] = 8'h8c;
    mem[12'h02b6] = 8'h15;
    mem[12'h02b7] = 8'h15;
    mem[12'h02b8] = 8'h08;
    mem[12'h02b9] = 8'h14;
    mem[12'h02ba] = 8'h38;
    mem[12'h02bb] = 8'h8c;
    mem[12'h02bc] = 8'h15;
    mem[12'h02bd] = 8'h15;
    mem[12'h02be] = 8'h08;
    mem[12'h02bf] = 8'h15;
    mem[12'h02c0] = 8'h37;
    mem[12'h02c1] = 8'h27;
    mem[12'h02c2] = 8'h15;
    mem[12'h02c3] = 8'h27;
    mem[12'h02c4] = 8'h3b;
    mem[12'h02c5] = 8'h15;
    mem[12'h02c6] = 8'h09;
    mem[12'h02c7] = 8'h15;
    mem[12'h02c8] = 8'h37;
    mem[12'h02c9] = 8'h27;
    mem[12'h02ca] = 8'h15;
    mem[12'h02cb] = 8'h27;
    mem[12'h02cc] = 8'h3b;
    mem[12'h02cd] = 8'h15;
    mem[12'h02ce] = 8'h09;
    mem[12'h02cf] = 8'h15;
    mem[12'h02d0] = 8'h37;
    mem[12'h02d1] = 8'h27;
    mem[12'h02d2] = 8'h15;
    mem[12'h02d3] = 8'h27;
    mem[12'h02d4] = 8'h3b;
    mem[12'h02d5] = 8'h15;
    mem[12'h02d6] = 8'h09;
    mem[12'h02d7] = 8'h15;
    mem[12'h02d8] = 8'h37;
    mem[12'h02d9] = 8'h27;
    mem[12'h02da] = 8'h15;
    mem[12'h02db] = 8'h27;
    mem[12'h02dc] = 8'h3b;
    mem[12'h02dd] = 8'h15;
    mem[12'h02de] = 8'h0a;
    mem[12'h02df] = 8'h15;
    mem[12'h02e0] = 8'h36;
    mem[12'h02e1] = 8'h27;
    mem[12'h02e2] = 8'h15;
    mem[12'h02e3] = 8'h27;
    mem[12'h02e4] = 8'h3a;
    mem[12'h02e5] = 8'h16;
    mem[12'h02e6] = 8'h0a;
    mem[12'h02e7] = 8'h15;
    mem[12'h02e8] = 8'h36;
    mem[12'h02e9] = 8'h27;
    mem[12'h02ea] = 8'h15;
    mem[12'h02eb] = 8'h27;
    mem[12'h02ec] = 8'h3a;
    mem[12'h02ed] = 8'h15;
    mem[12'h02ee] = 8'h0b;
    mem[12'h02ef] = 8'h15;
    mem[12'h02f0] = 8'h36;
    mem[12'h02f1] = 8'h27;
    mem[12'h02f2] = 8'h15;
    mem[12'h02f3] = 8'h27;
    mem[12'h02f4] = 8'h3a;
    mem[12'h02f5] = 8'h15;
    mem[12'h02f6] = 8'h0b;
    mem[12'h02f7] = 8'h16;
    mem[12'h02f8] = 8'h35;
    mem[12'h02f9] = 8'h27;
    mem[12'h02fa] = 8'h15;
    mem[12'h02fb] = 8'h27;
    mem[12'h02fc] = 8'h39;
    mem[12'h02fd] = 8'h16;
    mem[12'h02fe] = 8'h0c;
    mem[12'h02ff] = 8'h15;
    mem[12'h0300] = 8'h35;
    mem[12'h0301] = 8'h27;
    mem[12'h0302] = 8'h15;
    mem[12'h0303] = 8'h27;
    mem[12'h0304] = 8'h39;
    mem[12'h0305] = 8'h16;
    mem[12'h0306] = 8'h0c;
    mem[12'h0307] = 8'h15;
    mem[12'h0308] = 8'h35;
    mem[12'h0309] = 8'h27;
    mem[12'h030a] = 8'h15;
    mem[12'h030b] = 8'h27;
    mem[12'h030c] = 8'h39;
    mem[12'h030d] = 8'h15;
    mem[12'h030e] = 8'h0d;
    mem[12'h030f] = 8'h16;
    mem[12'h0310] = 8'h34;
    mem[12'h0311] = 8'h27;
    mem[12'h0312] = 8'h15;
    mem[12'h0313] = 8'h27;
    mem[12'h0314] = 8'h39;
    mem[12'h0315] = 8'h15;
    mem[12'h0316] = 8'h0d;
    mem[12'h0317] = 8'h16;
    mem[12'h0318] = 8'h34;
    mem[12'h0319] = 8'h27;
    mem[12'h031a] = 8'h15;
    mem[12'h031b] = 8'h27;
    mem[12'h031c] = 8'h38;
    mem[12'h031d] = 8'h16;
    mem[12'h031e] = 8'h0e;
    mem[12'h031f] = 8'h15;
    mem[12'h0320] = 8'h34;
    mem[12'h0321] = 8'h27;
    mem[12'h0322] = 8'h15;
    mem[12'h0323] = 8'h27;
    mem[12'h0324] = 8'h38;
    mem[12'h0325] = 8'h16;
    mem[12'h0326] = 8'h0e;
    mem[12'h0327] = 8'h16;
    mem[12'h0328] = 8'h33;
    mem[12'h0329] = 8'h27;
    mem[12'h032a] = 8'h15;
    mem[12'h032b] = 8'h27;
    mem[12'h032c] = 8'h37;
    mem[12'h032d] = 8'h16;
    mem[12'h032e] = 8'h0f;
    mem[12'h032f] = 8'h16;
    mem[12'h0330] = 8'h33;
    mem[12'h0331] = 8'h27;
    mem[12'h0332] = 8'h15;
    mem[12'h0333] = 8'h27;
    mem[12'h0334] = 8'h37;
    mem[12'h0335] = 8'h16;
    mem[12'h0336] = 8'h10;
    mem[12'h0337] = 8'h15;
    mem[12'h0338] = 8'h33;
    mem[12'h0339] = 8'h27;
    mem[12'h033a] = 8'h15;
    mem[12'h033b] = 8'h27;
    mem[12'h033c] = 8'h37;
    mem[12'h033d] = 8'h16;
    mem[12'h033e] = 8'h10;
    mem[12'h033f] = 8'h16;
    mem[12'h0340] = 8'h32;
    mem[12'h0341] = 8'h27;
    mem[12'h0342] = 8'h15;
    mem[12'h0343] = 8'h27;
    mem[12'h0344] = 8'h36;
    mem[12'h0345] = 8'h16;
    mem[12'h0346] = 8'h11;
    mem[12'h0347] = 8'h16;
    mem[12'h0348] = 8'h32;
    mem[12'h0349] = 8'h27;
    mem[12'h034a] = 8'h15;
    mem[12'h034b] = 8'h27;
    mem[12'h034c] = 8'h36;
    mem[12'h034d] = 8'h16;
    mem[12'h034e] = 8'h12;
    mem[12'h034f] = 8'h16;
    mem[12'h0350] = 8'h31;
    mem[12'h0351] = 8'h27;
    mem[12'h0352] = 8'h15;
    mem[12'h0353] = 8'h27;
    mem[12'h0354] = 8'h35;
    mem[12'h0355] = 8'h17;
    mem[12'h0356] = 8'h12;
    mem[12'h0357] = 8'h16;
    mem[12'h0358] = 8'h31;
    mem[12'h0359] = 8'h27;
    mem[12'h035a] = 8'h15;
    mem[12'h035b] = 8'h27;
    mem[12'h035c] = 8'h35;
    mem[12'h035d] = 8'h16;
    mem[12'h035e] = 8'h13;
    mem[12'h035f] = 8'h16;
    mem[12'h0360] = 8'h31;
    mem[12'h0361] = 8'h27;
    mem[12'h0362] = 8'h15;
    mem[12'h0363] = 8'h27;
    mem[12'h0364] = 8'h35;
    mem[12'h0365] = 8'h16;
    mem[12'h0366] = 8'h14;
    mem[12'h0367] = 8'h16;
    mem[12'h0368] = 8'h30;
    mem[12'h0369] = 8'h27;
    mem[12'h036a] = 8'h15;
    mem[12'h036b] = 8'h27;
    mem[12'h036c] = 8'h34;
    mem[12'h036d] = 8'h17;
    mem[12'h036e] = 8'h14;
    mem[12'h036f] = 8'h16;
    mem[12'h0370] = 8'h30;
    mem[12'h0371] = 8'h27;
    mem[12'h0372] = 8'h15;
    mem[12'h0373] = 8'h27;
    mem[12'h0374] = 8'h34;
    mem[12'h0375] = 8'h16;
    mem[12'h0376] = 8'h15;
    mem[12'h0377] = 8'h17;
    mem[12'h0378] = 8'h2f;
    mem[12'h0379] = 8'h27;
    mem[12'h037a] = 8'h15;
    mem[12'h037b] = 8'h27;
    mem[12'h037c] = 8'h33;
    mem[12'h037d] = 8'h17;
    mem[12'h037e] = 8'h16;
    mem[12'h037f] = 8'h16;
    mem[12'h0380] = 8'h6d;
    mem[12'h0381] = 8'h27;
    mem[12'h0382] = 8'h33;
    mem[12'h0383] = 8'h16;
    mem[12'h0384] = 8'h17;
    mem[12'h0385] = 8'h17;
    mem[12'h0386] = 8'h6c;
    mem[12'h0387] = 8'h27;
    mem[12'h0388] = 8'h32;
    mem[12'h0389] = 8'h17;
    mem[12'h038a] = 8'h18;
    mem[12'h038b] = 8'h16;
    mem[12'h038c] = 8'h6c;
    mem[12'h038d] = 8'h27;
    mem[12'h038e] = 8'h32;
    mem[12'h038f] = 8'h17;
    mem[12'h0390] = 8'h18;
    mem[12'h0391] = 8'h17;
    mem[12'h0392] = 8'h6b;
    mem[12'h0393] = 8'h27;
    mem[12'h0394] = 8'h31;
    mem[12'h0395] = 8'h17;
    mem[12'h0396] = 8'h19;
    mem[12'h0397] = 8'h17;
    mem[12'h0398] = 8'h6b;
    mem[12'h0399] = 8'h27;
    mem[12'h039a] = 8'h31;
    mem[12'h039b] = 8'h17;
    mem[12'h039c] = 8'h1a;
    mem[12'h039d] = 8'h17;
    mem[12'h039e] = 8'h6a;
    mem[12'h039f] = 8'h27;
    mem[12'h03a0] = 8'h30;
    mem[12'h03a1] = 8'h17;
    mem[12'h03a2] = 8'h1b;
    mem[12'h03a3] = 8'h18;
    mem[12'h03a4] = 8'h69;
    mem[12'h03a5] = 8'h27;
    mem[12'h03a6] = 8'h30;
    mem[12'h03a7] = 8'h17;
    mem[12'h03a8] = 8'h1c;
    mem[12'h03a9] = 8'h17;
    mem[12'h03aa] = 8'h69;
    mem[12'h03ab] = 8'h27;
    mem[12'h03ac] = 8'h2f;
    mem[12'h03ad] = 8'h17;
    mem[12'h03ae] = 8'h1d;
    mem[12'h03af] = 8'h18;
    mem[12'h03b0] = 8'h68;
    mem[12'h03b1] = 8'h27;
    mem[12'h03b2] = 8'h2e;
    mem[12'h03b3] = 8'h18;
    mem[12'h03b4] = 8'h1e;
    mem[12'h03b5] = 8'h17;
    mem[12'h03b6] = 8'h68;
    mem[12'h03b7] = 8'h27;
    mem[12'h03b8] = 8'h2e;
    mem[12'h03b9] = 8'h17;
    mem[12'h03ba] = 8'h1f;
    mem[12'h03bb] = 8'h18;
    mem[12'h03bc] = 8'h67;
    mem[12'h03bd] = 8'h27;
    mem[12'h03be] = 8'h2d;
    mem[12'h03bf] = 8'h18;
    mem[12'h03c0] = 8'h20;
    mem[12'h03c1] = 8'h18;
    mem[12'h03c2] = 8'h66;
    mem[12'h03c3] = 8'h27;
    mem[12'h03c4] = 8'h2d;
    mem[12'h03c5] = 8'h17;
    mem[12'h03c6] = 8'h21;
    mem[12'h03c7] = 8'h18;
    mem[12'h03c8] = 8'h66;
    mem[12'h03c9] = 8'h27;
    mem[12'h03ca] = 8'h2c;
    mem[12'h03cb] = 8'h18;
    mem[12'h03cc] = 8'h22;
    mem[12'h03cd] = 8'h18;
    mem[12'h03ce] = 8'h65;
    mem[12'h03cf] = 8'h27;
    mem[12'h03d0] = 8'h2b;
    mem[12'h03d1] = 8'h18;
    mem[12'h03d2] = 8'h23;
    mem[12'h03d3] = 8'h19;
    mem[12'h03d4] = 8'h64;
    mem[12'h03d5] = 8'h27;
    mem[12'h03d6] = 8'h2a;
    mem[12'h03d7] = 8'h19;
    mem[12'h03d8] = 8'h24;
    mem[12'h03d9] = 8'h18;
    mem[12'h03da] = 8'h64;
    mem[12'h03db] = 8'h27;
    mem[12'h03dc] = 8'h2a;
    mem[12'h03dd] = 8'h18;
    mem[12'h03de] = 8'h25;
    mem[12'h03df] = 8'h19;
    mem[12'h03e0] = 8'h63;
    mem[12'h03e1] = 8'h27;
    mem[12'h03e2] = 8'h29;
    mem[12'h03e3] = 8'h19;
    mem[12'h03e4] = 8'h26;
    mem[12'h03e5] = 8'h19;
    mem[12'h03e6] = 8'h62;
    mem[12'h03e7] = 8'h27;
    mem[12'h03e8] = 8'h28;
    mem[12'h03e9] = 8'h19;
    mem[12'h03ea] = 8'h28;
    mem[12'h03eb] = 8'h18;
    mem[12'h03ec] = 8'h62;
    mem[12'h03ed] = 8'h27;
    mem[12'h03ee] = 8'h28;
    mem[12'h03ef] = 8'h19;
    mem[12'h03f0] = 8'h28;
    mem[12'h03f1] = 8'h19;
    mem[12'h03f2] = 8'h61;
    mem[12'h03f3] = 8'h27;
    mem[12'h03f4] = 8'h27;
    mem[12'h03f5] = 8'h19;
    mem[12'h03f6] = 8'h2a;
    mem[12'h03f7] = 8'h19;
    mem[12'h03f8] = 8'h60;
    mem[12'h03f9] = 8'h27;
    mem[12'h03fa] = 8'h26;
    mem[12'h03fb] = 8'h19;
    mem[12'h03fc] = 8'h2b;
    mem[12'h03fd] = 8'h1a;
    mem[12'h03fe] = 8'h5f;
    mem[12'h03ff] = 8'h27;
    mem[12'h0400] = 8'h25;
    mem[12'h0401] = 8'h1a;
    mem[12'h0402] = 8'h2c;
    mem[12'h0403] = 8'h1a;
    mem[12'h0404] = 8'h5e;
    mem[12'h0405] = 8'h27;
    mem[12'h0406] = 8'h24;
    mem[12'h0407] = 8'h1a;
    mem[12'h0408] = 8'h2e;
    mem[12'h0409] = 8'h19;
    mem[12'h040a] = 8'h5e;
    mem[12'h040b] = 8'h27;
    mem[12'h040c] = 8'h24;
    mem[12'h040d] = 8'h1a;
    mem[12'h040e] = 8'h2e;
    mem[12'h040f] = 8'h1a;
    mem[12'h0410] = 8'h5d;
    mem[12'h0411] = 8'h27;
    mem[12'h0412] = 8'h23;
    mem[12'h0413] = 8'h1a;
    mem[12'h0414] = 8'h30;
    mem[12'h0415] = 8'h1a;
    mem[12'h0416] = 8'h5c;
    mem[12'h0417] = 8'h27;
    mem[12'h0418] = 8'h22;
    mem[12'h0419] = 8'h1a;
    mem[12'h041a] = 8'h32;
    mem[12'h041b] = 8'h1a;
    mem[12'h041c] = 8'h5b;
    mem[12'h041d] = 8'h27;
    mem[12'h041e] = 8'h21;
    mem[12'h041f] = 8'h1b;
    mem[12'h0420] = 8'h32;
    mem[12'h0421] = 8'h1b;
    mem[12'h0422] = 8'h5a;
    mem[12'h0423] = 8'h27;
    mem[12'h0424] = 8'h20;
    mem[12'h0425] = 8'h1b;
    mem[12'h0426] = 8'h34;
    mem[12'h0427] = 8'h1b;
    mem[12'h0428] = 8'h59;
    mem[12'h0429] = 8'h27;
    mem[12'h042a] = 8'h1f;
    mem[12'h042b] = 8'h1b;
    mem[12'h042c] = 8'h36;
    mem[12'h042d] = 8'h1b;
    mem[12'h042e] = 8'h58;
    mem[12'h042f] = 8'h27;
    mem[12'h0430] = 8'h1e;
    mem[12'h0431] = 8'h1b;
    mem[12'h0432] = 8'h37;
    mem[12'h0433] = 8'h1c;
    mem[12'h0434] = 8'h57;
    mem[12'h0435] = 8'h27;
    mem[12'h0436] = 8'h1d;
    mem[12'h0437] = 8'h1c;
    mem[12'h0438] = 8'h38;
    mem[12'h0439] = 8'h1c;
    mem[12'h043a] = 8'h56;
    mem[12'h043b] = 8'h27;
    mem[12'h043c] = 8'h1c;
    mem[12'h043d] = 8'h1c;
    mem[12'h043e] = 8'h3a;
    mem[12'h043f] = 8'h1c;
    mem[12'h0440] = 8'h55;
    mem[12'h0441] = 8'h27;
    mem[12'h0442] = 8'h1b;
    mem[12'h0443] = 8'h1c;
    mem[12'h0444] = 8'h3c;
    mem[12'h0445] = 8'h1c;
    mem[12'h0446] = 8'h54;
    mem[12'h0447] = 8'h27;
    mem[12'h0448] = 8'h1a;
    mem[12'h0449] = 8'h1c;
    mem[12'h044a] = 8'h3e;
    mem[12'h044b] = 8'h1c;
    mem[12'h044c] = 8'h53;
    mem[12'h044d] = 8'h27;
    mem[12'h044e] = 8'h19;
    mem[12'h044f] = 8'h1d;
    mem[12'h0450] = 8'h3e;
    mem[12'h0451] = 8'h1d;
    mem[12'h0452] = 8'h52;
    mem[12'h0453] = 8'h27;
    mem[12'h0454] = 8'h18;
    mem[12'h0455] = 8'h1d;
    mem[12'h0456] = 8'h40;
    mem[12'h0457] = 8'h1d;
    mem[12'h0458] = 8'h51;
    mem[12'h0459] = 8'h27;
    mem[12'h045a] = 8'h17;
    mem[12'h045b] = 8'h1d;
    mem[12'h045c] = 8'h42;
    mem[12'h045d] = 8'h1e;
    mem[12'h045e] = 8'h4f;
    mem[12'h045f] = 8'h27;
    mem[12'h0460] = 8'h15;
    mem[12'h0461] = 8'h1e;
    mem[12'h0462] = 8'h44;
    mem[12'h0463] = 8'h1e;
    mem[12'h0464] = 8'h4e;
    mem[12'h0465] = 8'h27;
    mem[12'h0466] = 8'h14;
    mem[12'h0467] = 8'h1e;
    mem[12'h0468] = 8'h46;
    mem[12'h0469] = 8'h1e;
    mem[12'h046a] = 8'h4d;
    mem[12'h046b] = 8'h27;
    mem[12'h046c] = 8'h13;
    mem[12'h046d] = 8'h1e;
    mem[12'h046e] = 8'h48;
    mem[12'h046f] = 8'h1e;
    mem[12'h0470] = 8'h4c;
    mem[12'h0471] = 8'h27;
    mem[12'h0472] = 8'h12;
    mem[12'h0473] = 8'h1e;
    mem[12'h0474] = 8'h49;
    mem[12'h0475] = 8'h20;
    mem[12'h0476] = 8'h4a;
    mem[12'h0477] = 8'h27;
    mem[12'h0478] = 8'h10;
    mem[12'h0479] = 8'h20;
    mem[12'h047a] = 8'h4a;
    mem[12'h047b] = 8'h20;
    mem[12'h047c] = 8'h49;
    mem[12'h047d] = 8'h27;
    mem[12'h047e] = 8'h0f;
    mem[12'h047f] = 8'h20;
    mem[12'h0480] = 8'h4c;
    mem[12'h0481] = 8'h21;
    mem[12'h0482] = 8'h47;
    mem[12'h0483] = 8'h27;
    mem[12'h0484] = 8'h0d;
    mem[12'h0485] = 8'h21;
    mem[12'h0486] = 8'h4e;
    mem[12'h0487] = 8'h21;
    mem[12'h0488] = 8'h46;
    mem[12'h0489] = 8'h27;
    mem[12'h048a] = 8'h0c;
    mem[12'h048b] = 8'h21;
    mem[12'h048c] = 8'h50;
    mem[12'h048d] = 8'h22;
    mem[12'h048e] = 8'h44;
    mem[12'h048f] = 8'h27;
    mem[12'h0490] = 8'h0b;
    mem[12'h0491] = 8'h21;
    mem[12'h0492] = 8'h52;
    mem[12'h0493] = 8'h22;
    mem[12'h0494] = 8'h43;
    mem[12'h0495] = 8'h27;
    mem[12'h0496] = 8'h0a;
    mem[12'h0497] = 8'h21;
    mem[12'h0498] = 8'h54;
    mem[12'h0499] = 8'h23;
    mem[12'h049a] = 8'h41;
    mem[12'h049b] = 8'h27;
    mem[12'h049c] = 8'h0a;
    mem[12'h049d] = 8'h20;
    mem[12'h049e] = 8'h56;
    mem[12'h049f] = 8'h24;
    mem[12'h04a0] = 8'h3f;
    mem[12'h04a1] = 8'h27;
    mem[12'h04a2] = 8'h0a;
    mem[12'h04a3] = 8'h1f;
    mem[12'h04a4] = 8'h58;
    mem[12'h04a5] = 8'h24;
    mem[12'h04a6] = 8'h3e;
    mem[12'h04a7] = 8'h27;
    mem[12'h04a8] = 8'h0a;
    mem[12'h04a9] = 8'h1e;
    mem[12'h04aa] = 8'h5b;
    mem[12'h04ab] = 8'h24;
    mem[12'h04ac] = 8'h3c;
    mem[12'h04ad] = 8'h27;
    mem[12'h04ae] = 8'h0a;
    mem[12'h04af] = 8'h1d;
    mem[12'h04b0] = 8'h5d;
    mem[12'h04b1] = 8'h25;
    mem[12'h04b2] = 8'h3a;
    mem[12'h04b3] = 8'h27;
    mem[12'h04b4] = 8'h0a;
    mem[12'h04b5] = 8'h1b;
    mem[12'h04b6] = 8'h60;
    mem[12'h04b7] = 8'h26;
    mem[12'h04b8] = 8'h38;
    mem[12'h04b9] = 8'h27;
    mem[12'h04ba] = 8'h0a;
    mem[12'h04bb] = 8'h1a;
    mem[12'h04bc] = 8'h62;
    mem[12'h04bd] = 8'h27;
    mem[12'h04be] = 8'h36;
    mem[12'h04bf] = 8'h27;
    mem[12'h04c0] = 8'h0a;
    mem[12'h04c1] = 8'h19;
    mem[12'h04c2] = 8'h64;
    mem[12'h04c3] = 8'h29;
    mem[12'h04c4] = 8'h33;
    mem[12'h04c5] = 8'h27;
    mem[12'h04c6] = 8'h0a;
    mem[12'h04c7] = 8'h18;
    mem[12'h04c8] = 8'h67;
    mem[12'h04c9] = 8'h29;
    mem[12'h04ca] = 8'h31;
    mem[12'h04cb] = 8'h27;
    mem[12'h04cc] = 8'h0a;
    mem[12'h04cd] = 8'h17;
    mem[12'h04ce] = 8'h69;
    mem[12'h04cf] = 8'h2b;
    mem[12'h04d0] = 8'h2e;
    mem[12'h04d1] = 8'h27;
    mem[12'h04d2] = 8'h0a;
    mem[12'h04d3] = 8'h15;
    mem[12'h04d4] = 8'h6c;
    mem[12'h04d5] = 8'h2d;
    mem[12'h04d6] = 8'h2b;
    mem[12'h04d7] = 8'h27;
    mem[12'h04d8] = 8'h0a;
    mem[12'h04d9] = 8'h14;
    mem[12'h04da] = 8'h6e;
    mem[12'h04db] = 8'h2f;
    mem[12'h04dc] = 8'h28;
    mem[12'h04dd] = 8'h27;
    mem[12'h04de] = 8'h0a;
    mem[12'h04df] = 8'h13;
    mem[12'h04e0] = 8'h71;
    mem[12'h04e1] = 8'h30;
    mem[12'h04e2] = 8'h25;
    mem[12'h04e3] = 8'h27;
    mem[12'h04e4] = 8'h0a;
    mem[12'h04e5] = 8'h11;
    mem[12'h04e6] = 8'h74;
    mem[12'h04e7] = 8'h33;
    mem[12'h04e8] = 8'h21;
    mem[12'h04e9] = 8'h27;
    mem[12'h04ea] = 8'h0a;
    mem[12'h04eb] = 8'h10;
    mem[12'h04ec] = 8'h77;
    mem[12'h04ed] = 8'h36;
    mem[12'h04ee] = 8'h1c;
    mem[12'h04ef] = 8'h27;
    mem[12'h04f0] = 8'h0a;
    mem[12'h04f1] = 8'h0f;
    mem[12'h04f2] = 8'h79;
    mem[12'h04f3] = 8'h3c;
    mem[12'h04f4] = 8'h15;
    mem[12'h04f5] = 8'h27;
    mem[12'h04f6] = 8'h0a;
    mem[12'h04f7] = 8'h0d;
    mem[12'h04f8] = 8'h7d;
    mem[12'h04f9] = 8'h78;
    mem[12'h04fa] = 8'h0a;
    mem[12'h04fb] = 8'h0c;
    mem[12'h04fc] = 8'h7f;
    mem[12'h04fd] = 8'h77;
    mem[12'h04fe] = 8'h0a;
    mem[12'h04ff] = 8'h0a;
    mem[12'h0500] = 8'h83;
    mem[12'h0501] = 8'h75;
    mem[12'h0502] = 8'h0a;
    mem[12'h0503] = 8'h08;
    mem[12'h0504] = 8'h87;
    mem[12'h0505] = 8'h73;
    mem[12'h0506] = 8'h0a;
    mem[12'h0507] = 8'h07;
    mem[12'h0508] = 8'h89;
    mem[12'h0509] = 8'h72;
    mem[12'h050a] = 8'h0a;
    mem[12'h050b] = 8'h05;
    mem[12'h050c] = 8'h8d;
    mem[12'h050d] = 8'h70;
    mem[12'h050e] = 8'h0a;
    mem[12'h050f] = 8'h03;
    mem[12'h0510] = 8'h91;
    mem[12'h0511] = 8'h6e;
    mem[12'h0512] = 8'h0a;
    mem[12'h0513] = 8'h01;
    mem[12'h0514] = 8'h95;
    mem[12'h0515] = 8'h6c;
    mem[12'h0516] = 8'ha4;
    mem[12'h0517] = 8'h6a;
    mem[12'h0518] = 8'ha6;
    mem[12'h0519] = 8'h68;
    mem[12'h051a] = 8'ha8;
    mem[12'h051b] = 8'h66;
    mem[12'h051c] = 8'hab;
    mem[12'h051d] = 8'h63;
    mem[12'h051e] = 8'had;
    mem[12'h051f] = 8'h61;
    mem[12'h0520] = 8'hb0;
    mem[12'h0521] = 8'h5b;
    mem[12'h0522] = 8'hb6;
    mem[12'h0523] = 8'h55;
    mem[12'h0524] = 8'hbc;
    mem[12'h0525] = 8'h4f;
    mem[12'h0526] = 8'hc2;
    mem[12'h0527] = 8'h49;
    mem[12'h0528] = 8'hc9;
    mem[12'h0529] = 8'h41;
    mem[12'h052a] = 8'hd1;
    mem[12'h052b] = 8'h39;
    mem[12'h052c] = 8'hda;
    mem[12'h052d] = 8'h2f;
    mem[12'h052e] = 8'he5;
    mem[12'h052f] = 8'h22;
    mem[12'h0530] = 8'hf9;
    mem[12'h0531] = 8'h0a;
  end
  assign len = mem[addr];
endmodule



module bitmap_rom (
    input wire [6:0] x,
    input wire [6:0] y,
    output wire pixel
);

  reg [7:0] mem[2047:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h80;
    mem[23] = 8'hff;
    mem[24] = 8'hff;
    mem[25] = 8'h01;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'hfc;
    mem[39] = 8'hff;
    mem[40] = 8'hff;
    mem[41] = 8'h3f;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'hc0;
    mem[54] = 8'hff;
    mem[55] = 8'hff;
    mem[56] = 8'hff;
    mem[57] = 8'hff;
    mem[58] = 8'h03;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'hf8;
    mem[70] = 8'hff;
    mem[71] = 8'hff;
    mem[72] = 8'hff;
    mem[73] = 8'hff;
    mem[74] = 8'h1f;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'hff;
    mem[86] = 8'hff;
    mem[87] = 8'hff;
    mem[88] = 8'hff;
    mem[89] = 8'hff;
    mem[90] = 8'hff;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'hc0;
    mem[101] = 8'hff;
    mem[102] = 8'hff;
    mem[103] = 8'hff;
    mem[104] = 8'hff;
    mem[105] = 8'hff;
    mem[106] = 8'hff;
    mem[107] = 8'h03;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'hf0;
    mem[117] = 8'hff;
    mem[118] = 8'hff;
    mem[119] = 8'hff;
    mem[120] = 8'hff;
    mem[121] = 8'hff;
    mem[122] = 8'hff;
    mem[123] = 8'h0f;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'hfc;
    mem[133] = 8'hff;
    mem[134] = 8'hff;
    mem[135] = 8'hff;
    mem[136] = 8'hff;
    mem[137] = 8'hff;
    mem[138] = 8'hff;
    mem[139] = 8'h3f;
    mem[140] = 8'h00;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'hff;
    mem[149] = 8'hff;
    mem[150] = 8'hff;
    mem[151] = 8'hff;
    mem[152] = 8'hff;
    mem[153] = 8'hff;
    mem[154] = 8'hff;
    mem[155] = 8'hff;
    mem[156] = 8'h00;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h00;
    mem[162] = 8'h00;
    mem[163] = 8'hc0;
    mem[164] = 8'hff;
    mem[165] = 8'hff;
    mem[166] = 8'hff;
    mem[167] = 8'hff;
    mem[168] = 8'hff;
    mem[169] = 8'hff;
    mem[170] = 8'hff;
    mem[171] = 8'hff;
    mem[172] = 8'h03;
    mem[173] = 8'h00;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h00;
    mem[178] = 8'h00;
    mem[179] = 8'he0;
    mem[180] = 8'hff;
    mem[181] = 8'hff;
    mem[182] = 8'hff;
    mem[183] = 8'h7f;
    mem[184] = 8'hfe;
    mem[185] = 8'hff;
    mem[186] = 8'hff;
    mem[187] = 8'hff;
    mem[188] = 8'h07;
    mem[189] = 8'h00;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
    mem[192] = 8'h00;
    mem[193] = 8'h00;
    mem[194] = 8'h00;
    mem[195] = 8'hf8;
    mem[196] = 8'hff;
    mem[197] = 8'hff;
    mem[198] = 8'h3f;
    mem[199] = 8'h00;
    mem[200] = 8'h00;
    mem[201] = 8'hfc;
    mem[202] = 8'hff;
    mem[203] = 8'hff;
    mem[204] = 8'h1f;
    mem[205] = 8'h00;
    mem[206] = 8'h00;
    mem[207] = 8'h00;
    mem[208] = 8'h00;
    mem[209] = 8'h00;
    mem[210] = 8'h00;
    mem[211] = 8'hfc;
    mem[212] = 8'hff;
    mem[213] = 8'hff;
    mem[214] = 8'h03;
    mem[215] = 8'h00;
    mem[216] = 8'h00;
    mem[217] = 8'hc0;
    mem[218] = 8'hff;
    mem[219] = 8'hff;
    mem[220] = 8'h3f;
    mem[221] = 8'h00;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'h00;
    mem[227] = 8'hfe;
    mem[228] = 8'hff;
    mem[229] = 8'h7f;
    mem[230] = 8'h00;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'hfe;
    mem[235] = 8'hff;
    mem[236] = 8'h7f;
    mem[237] = 8'h00;
    mem[238] = 8'h00;
    mem[239] = 8'h00;
    mem[240] = 8'h00;
    mem[241] = 8'h00;
    mem[242] = 8'h80;
    mem[243] = 8'hff;
    mem[244] = 8'hff;
    mem[245] = 8'h0f;
    mem[246] = 8'h00;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'hf0;
    mem[251] = 8'hff;
    mem[252] = 8'hff;
    mem[253] = 8'h01;
    mem[254] = 8'h00;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'h00;
    mem[258] = 8'hc0;
    mem[259] = 8'hff;
    mem[260] = 8'hff;
    mem[261] = 8'h03;
    mem[262] = 8'h00;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'hc0;
    mem[267] = 8'hff;
    mem[268] = 8'hff;
    mem[269] = 8'h03;
    mem[270] = 8'h00;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'he0;
    mem[275] = 8'hff;
    mem[276] = 8'hff;
    mem[277] = 8'h00;
    mem[278] = 8'h00;
    mem[279] = 8'h00;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'h00;
    mem[283] = 8'hff;
    mem[284] = 8'hff;
    mem[285] = 8'h07;
    mem[286] = 8'h00;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'hf0;
    mem[291] = 8'hff;
    mem[292] = 8'h3f;
    mem[293] = 8'h00;
    mem[294] = 8'h00;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'h00;
    mem[299] = 8'hfc;
    mem[300] = 8'hff;
    mem[301] = 8'h0f;
    mem[302] = 8'h00;
    mem[303] = 8'h00;
    mem[304] = 8'h00;
    mem[305] = 8'h00;
    mem[306] = 8'hf8;
    mem[307] = 8'hff;
    mem[308] = 8'h0f;
    mem[309] = 8'h00;
    mem[310] = 8'h00;
    mem[311] = 8'h00;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'h00;
    mem[315] = 8'hf0;
    mem[316] = 8'hff;
    mem[317] = 8'h1f;
    mem[318] = 8'h00;
    mem[319] = 8'h00;
    mem[320] = 8'h00;
    mem[321] = 8'h00;
    mem[322] = 8'hfc;
    mem[323] = 8'hff;
    mem[324] = 8'h07;
    mem[325] = 8'h00;
    mem[326] = 8'h00;
    mem[327] = 8'h00;
    mem[328] = 8'h00;
    mem[329] = 8'h00;
    mem[330] = 8'h00;
    mem[331] = 8'he0;
    mem[332] = 8'hff;
    mem[333] = 8'h3f;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
    mem[336] = 8'h00;
    mem[337] = 8'h00;
    mem[338] = 8'hfe;
    mem[339] = 8'hff;
    mem[340] = 8'h01;
    mem[341] = 8'h00;
    mem[342] = 8'h00;
    mem[343] = 8'h00;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'h00;
    mem[347] = 8'h80;
    mem[348] = 8'hff;
    mem[349] = 8'h7f;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'h00;
    mem[354] = 8'hff;
    mem[355] = 8'hff;
    mem[356] = 8'h00;
    mem[357] = 8'h00;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'hff;
    mem[365] = 8'hff;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h80;
    mem[370] = 8'hff;
    mem[371] = 8'h7f;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'hfe;
    mem[381] = 8'hff;
    mem[382] = 8'h01;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h80;
    mem[386] = 8'hff;
    mem[387] = 8'h3f;
    mem[388] = 8'h00;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'hfc;
    mem[397] = 8'hff;
    mem[398] = 8'h01;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'hc0;
    mem[402] = 8'hff;
    mem[403] = 8'h1f;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'hf8;
    mem[413] = 8'hff;
    mem[414] = 8'h03;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'he0;
    mem[418] = 8'hff;
    mem[419] = 8'h0f;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'he0;
    mem[429] = 8'hff;
    mem[430] = 8'h07;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'hf0;
    mem[434] = 8'hff;
    mem[435] = 8'hff;
    mem[436] = 8'hff;
    mem[437] = 8'hff;
    mem[438] = 8'hff;
    mem[439] = 8'hff;
    mem[440] = 8'hff;
    mem[441] = 8'h0f;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'hc0;
    mem[445] = 8'hff;
    mem[446] = 8'h0f;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'hf0;
    mem[450] = 8'hff;
    mem[451] = 8'hff;
    mem[452] = 8'hff;
    mem[453] = 8'hff;
    mem[454] = 8'hff;
    mem[455] = 8'hff;
    mem[456] = 8'hff;
    mem[457] = 8'h0f;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'hc0;
    mem[461] = 8'hff;
    mem[462] = 8'h0f;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'hf8;
    mem[466] = 8'hff;
    mem[467] = 8'hff;
    mem[468] = 8'hff;
    mem[469] = 8'hff;
    mem[470] = 8'hff;
    mem[471] = 8'hff;
    mem[472] = 8'hff;
    mem[473] = 8'h0f;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h80;
    mem[477] = 8'hff;
    mem[478] = 8'h1f;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'hfc;
    mem[482] = 8'hff;
    mem[483] = 8'hff;
    mem[484] = 8'hff;
    mem[485] = 8'hff;
    mem[486] = 8'hff;
    mem[487] = 8'hff;
    mem[488] = 8'hff;
    mem[489] = 8'h0f;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'hff;
    mem[494] = 8'h3f;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'hfc;
    mem[498] = 8'hff;
    mem[499] = 8'hff;
    mem[500] = 8'hff;
    mem[501] = 8'hff;
    mem[502] = 8'hff;
    mem[503] = 8'hff;
    mem[504] = 8'hff;
    mem[505] = 8'h0f;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'hfe;
    mem[510] = 8'h3f;
    mem[511] = 8'h00;
    mem[512] = 8'h00;
    mem[513] = 8'hfe;
    mem[514] = 8'hff;
    mem[515] = 8'hff;
    mem[516] = 8'hff;
    mem[517] = 8'hff;
    mem[518] = 8'hff;
    mem[519] = 8'hff;
    mem[520] = 8'hff;
    mem[521] = 8'h0f;
    mem[522] = 8'h00;
    mem[523] = 8'h00;
    mem[524] = 8'h00;
    mem[525] = 8'hfc;
    mem[526] = 8'h7f;
    mem[527] = 8'h00;
    mem[528] = 8'h00;
    mem[529] = 8'hfe;
    mem[530] = 8'hff;
    mem[531] = 8'hff;
    mem[532] = 8'hff;
    mem[533] = 8'hff;
    mem[534] = 8'hff;
    mem[535] = 8'hff;
    mem[536] = 8'hff;
    mem[537] = 8'h0f;
    mem[538] = 8'h00;
    mem[539] = 8'h00;
    mem[540] = 8'h00;
    mem[541] = 8'hf8;
    mem[542] = 8'h7f;
    mem[543] = 8'h00;
    mem[544] = 8'h00;
    mem[545] = 8'hff;
    mem[546] = 8'hff;
    mem[547] = 8'hff;
    mem[548] = 8'hff;
    mem[549] = 8'hff;
    mem[550] = 8'hff;
    mem[551] = 8'hff;
    mem[552] = 8'hff;
    mem[553] = 8'h0f;
    mem[554] = 8'h00;
    mem[555] = 8'h00;
    mem[556] = 8'h00;
    mem[557] = 8'hf8;
    mem[558] = 8'hff;
    mem[559] = 8'h00;
    mem[560] = 8'h00;
    mem[561] = 8'hff;
    mem[562] = 8'hff;
    mem[563] = 8'hff;
    mem[564] = 8'hff;
    mem[565] = 8'hff;
    mem[566] = 8'hff;
    mem[567] = 8'hff;
    mem[568] = 8'hff;
    mem[569] = 8'h0f;
    mem[570] = 8'h00;
    mem[571] = 8'h00;
    mem[572] = 8'h00;
    mem[573] = 8'hf0;
    mem[574] = 8'hff;
    mem[575] = 8'h00;
    mem[576] = 8'h80;
    mem[577] = 8'hff;
    mem[578] = 8'hff;
    mem[579] = 8'hff;
    mem[580] = 8'hff;
    mem[581] = 8'hff;
    mem[582] = 8'hff;
    mem[583] = 8'hff;
    mem[584] = 8'hff;
    mem[585] = 8'h0f;
    mem[586] = 8'h00;
    mem[587] = 8'h00;
    mem[588] = 8'h00;
    mem[589] = 8'he0;
    mem[590] = 8'hff;
    mem[591] = 8'h01;
    mem[592] = 8'h80;
    mem[593] = 8'hff;
    mem[594] = 8'hff;
    mem[595] = 8'hff;
    mem[596] = 8'hff;
    mem[597] = 8'hff;
    mem[598] = 8'hff;
    mem[599] = 8'hff;
    mem[600] = 8'hff;
    mem[601] = 8'h0f;
    mem[602] = 8'h00;
    mem[603] = 8'h00;
    mem[604] = 8'h00;
    mem[605] = 8'he0;
    mem[606] = 8'hff;
    mem[607] = 8'h01;
    mem[608] = 8'hc0;
    mem[609] = 8'hff;
    mem[610] = 8'hff;
    mem[611] = 8'hff;
    mem[612] = 8'hff;
    mem[613] = 8'hff;
    mem[614] = 8'hff;
    mem[615] = 8'hff;
    mem[616] = 8'hff;
    mem[617] = 8'h0f;
    mem[618] = 8'h00;
    mem[619] = 8'h00;
    mem[620] = 8'h00;
    mem[621] = 8'hc0;
    mem[622] = 8'hff;
    mem[623] = 8'h03;
    mem[624] = 8'hc0;
    mem[625] = 8'hff;
    mem[626] = 8'hff;
    mem[627] = 8'hff;
    mem[628] = 8'hff;
    mem[629] = 8'hff;
    mem[630] = 8'hff;
    mem[631] = 8'hff;
    mem[632] = 8'hff;
    mem[633] = 8'h0f;
    mem[634] = 8'h00;
    mem[635] = 8'h00;
    mem[636] = 8'h00;
    mem[637] = 8'hc0;
    mem[638] = 8'hff;
    mem[639] = 8'h03;
    mem[640] = 8'he0;
    mem[641] = 8'hff;
    mem[642] = 8'hff;
    mem[643] = 8'hff;
    mem[644] = 8'hff;
    mem[645] = 8'hff;
    mem[646] = 8'hff;
    mem[647] = 8'hff;
    mem[648] = 8'hff;
    mem[649] = 8'h0f;
    mem[650] = 8'h00;
    mem[651] = 8'h00;
    mem[652] = 8'h00;
    mem[653] = 8'h80;
    mem[654] = 8'hff;
    mem[655] = 8'h07;
    mem[656] = 8'he0;
    mem[657] = 8'hff;
    mem[658] = 8'hff;
    mem[659] = 8'hff;
    mem[660] = 8'hff;
    mem[661] = 8'hff;
    mem[662] = 8'hff;
    mem[663] = 8'hff;
    mem[664] = 8'hff;
    mem[665] = 8'h0f;
    mem[666] = 8'h00;
    mem[667] = 8'h00;
    mem[668] = 8'h00;
    mem[669] = 8'h80;
    mem[670] = 8'hff;
    mem[671] = 8'h07;
    mem[672] = 8'he0;
    mem[673] = 8'hff;
    mem[674] = 8'hff;
    mem[675] = 8'hff;
    mem[676] = 8'hff;
    mem[677] = 8'hff;
    mem[678] = 8'hff;
    mem[679] = 8'hff;
    mem[680] = 8'hff;
    mem[681] = 8'h0f;
    mem[682] = 8'h00;
    mem[683] = 8'h00;
    mem[684] = 8'h00;
    mem[685] = 8'h00;
    mem[686] = 8'hff;
    mem[687] = 8'h07;
    mem[688] = 8'hf0;
    mem[689] = 8'hff;
    mem[690] = 8'hff;
    mem[691] = 8'hff;
    mem[692] = 8'hff;
    mem[693] = 8'hff;
    mem[694] = 8'hff;
    mem[695] = 8'hff;
    mem[696] = 8'hff;
    mem[697] = 8'h0f;
    mem[698] = 8'h00;
    mem[699] = 8'h00;
    mem[700] = 8'h00;
    mem[701] = 8'h00;
    mem[702] = 8'hff;
    mem[703] = 8'h0f;
    mem[704] = 8'hf0;
    mem[705] = 8'hff;
    mem[706] = 8'hff;
    mem[707] = 8'hff;
    mem[708] = 8'hff;
    mem[709] = 8'hff;
    mem[710] = 8'hff;
    mem[711] = 8'hff;
    mem[712] = 8'hff;
    mem[713] = 8'h0f;
    mem[714] = 8'h00;
    mem[715] = 8'h00;
    mem[716] = 8'h00;
    mem[717] = 8'h00;
    mem[718] = 8'hfe;
    mem[719] = 8'h0f;
    mem[720] = 8'h00;
    mem[721] = 8'h00;
    mem[722] = 8'h00;
    mem[723] = 8'h00;
    mem[724] = 8'h80;
    mem[725] = 8'hff;
    mem[726] = 8'hff;
    mem[727] = 8'h03;
    mem[728] = 8'h00;
    mem[729] = 8'h00;
    mem[730] = 8'h00;
    mem[731] = 8'h00;
    mem[732] = 8'h00;
    mem[733] = 8'h00;
    mem[734] = 8'hfe;
    mem[735] = 8'h0f;
    mem[736] = 8'h00;
    mem[737] = 8'h00;
    mem[738] = 8'h00;
    mem[739] = 8'h00;
    mem[740] = 8'h80;
    mem[741] = 8'hff;
    mem[742] = 8'hff;
    mem[743] = 8'h03;
    mem[744] = 8'h00;
    mem[745] = 8'h00;
    mem[746] = 8'h00;
    mem[747] = 8'h00;
    mem[748] = 8'h00;
    mem[749] = 8'h00;
    mem[750] = 8'hfe;
    mem[751] = 8'h1f;
    mem[752] = 8'h00;
    mem[753] = 8'h00;
    mem[754] = 8'h00;
    mem[755] = 8'h00;
    mem[756] = 8'h80;
    mem[757] = 8'hff;
    mem[758] = 8'hff;
    mem[759] = 8'h03;
    mem[760] = 8'h00;
    mem[761] = 8'h00;
    mem[762] = 8'h00;
    mem[763] = 8'h00;
    mem[764] = 8'h00;
    mem[765] = 8'h00;
    mem[766] = 8'hfc;
    mem[767] = 8'h1f;
    mem[768] = 8'h00;
    mem[769] = 8'h00;
    mem[770] = 8'h00;
    mem[771] = 8'h00;
    mem[772] = 8'h80;
    mem[773] = 8'hff;
    mem[774] = 8'hff;
    mem[775] = 8'h03;
    mem[776] = 8'h00;
    mem[777] = 8'h00;
    mem[778] = 8'h00;
    mem[779] = 8'h00;
    mem[780] = 8'h00;
    mem[781] = 8'h00;
    mem[782] = 8'hfc;
    mem[783] = 8'h1f;
    mem[784] = 8'h00;
    mem[785] = 8'h00;
    mem[786] = 8'h00;
    mem[787] = 8'h00;
    mem[788] = 8'h80;
    mem[789] = 8'hff;
    mem[790] = 8'hff;
    mem[791] = 8'h03;
    mem[792] = 8'h00;
    mem[793] = 8'h00;
    mem[794] = 8'h00;
    mem[795] = 8'h00;
    mem[796] = 8'h00;
    mem[797] = 8'h00;
    mem[798] = 8'hfc;
    mem[799] = 8'h3f;
    mem[800] = 8'hfc;
    mem[801] = 8'h1f;
    mem[802] = 8'h00;
    mem[803] = 8'h00;
    mem[804] = 8'h80;
    mem[805] = 8'hff;
    mem[806] = 8'hff;
    mem[807] = 8'h03;
    mem[808] = 8'h00;
    mem[809] = 8'h00;
    mem[810] = 8'h00;
    mem[811] = 8'h00;
    mem[812] = 8'h00;
    mem[813] = 8'h00;
    mem[814] = 8'hf8;
    mem[815] = 8'h3f;
    mem[816] = 8'hfc;
    mem[817] = 8'h1f;
    mem[818] = 8'h00;
    mem[819] = 8'h00;
    mem[820] = 8'h80;
    mem[821] = 8'hff;
    mem[822] = 8'hff;
    mem[823] = 8'h03;
    mem[824] = 8'h00;
    mem[825] = 8'h00;
    mem[826] = 8'h00;
    mem[827] = 8'h00;
    mem[828] = 8'h00;
    mem[829] = 8'h00;
    mem[830] = 8'hf8;
    mem[831] = 8'h3f;
    mem[832] = 8'hfc;
    mem[833] = 8'h1f;
    mem[834] = 8'h00;
    mem[835] = 8'h00;
    mem[836] = 8'h80;
    mem[837] = 8'hff;
    mem[838] = 8'hff;
    mem[839] = 8'h03;
    mem[840] = 8'h00;
    mem[841] = 8'h00;
    mem[842] = 8'h00;
    mem[843] = 8'h00;
    mem[844] = 8'h00;
    mem[845] = 8'h00;
    mem[846] = 8'hf8;
    mem[847] = 8'h3f;
    mem[848] = 8'hfc;
    mem[849] = 8'h1f;
    mem[850] = 8'h00;
    mem[851] = 8'h00;
    mem[852] = 8'h80;
    mem[853] = 8'hff;
    mem[854] = 8'hff;
    mem[855] = 8'h03;
    mem[856] = 8'h00;
    mem[857] = 8'h00;
    mem[858] = 8'h00;
    mem[859] = 8'h00;
    mem[860] = 8'h00;
    mem[861] = 8'h00;
    mem[862] = 8'hf8;
    mem[863] = 8'h3f;
    mem[864] = 8'hfc;
    mem[865] = 8'h0f;
    mem[866] = 8'h00;
    mem[867] = 8'h00;
    mem[868] = 8'h80;
    mem[869] = 8'hff;
    mem[870] = 8'hff;
    mem[871] = 8'h03;
    mem[872] = 8'h00;
    mem[873] = 8'h00;
    mem[874] = 8'h00;
    mem[875] = 8'h00;
    mem[876] = 8'h00;
    mem[877] = 8'h00;
    mem[878] = 8'hf0;
    mem[879] = 8'h3f;
    mem[880] = 8'hfe;
    mem[881] = 8'h0f;
    mem[882] = 8'h00;
    mem[883] = 8'h00;
    mem[884] = 8'h80;
    mem[885] = 8'hff;
    mem[886] = 8'hff;
    mem[887] = 8'h03;
    mem[888] = 8'h00;
    mem[889] = 8'h00;
    mem[890] = 8'h00;
    mem[891] = 8'h00;
    mem[892] = 8'h00;
    mem[893] = 8'h00;
    mem[894] = 8'hf0;
    mem[895] = 8'h7f;
    mem[896] = 8'hfe;
    mem[897] = 8'h0f;
    mem[898] = 8'h00;
    mem[899] = 8'h00;
    mem[900] = 8'h80;
    mem[901] = 8'hff;
    mem[902] = 8'hff;
    mem[903] = 8'h03;
    mem[904] = 8'h00;
    mem[905] = 8'h00;
    mem[906] = 8'h00;
    mem[907] = 8'h00;
    mem[908] = 8'h00;
    mem[909] = 8'h00;
    mem[910] = 8'hf0;
    mem[911] = 8'h7f;
    mem[912] = 8'hfe;
    mem[913] = 8'h0f;
    mem[914] = 8'h00;
    mem[915] = 8'h00;
    mem[916] = 8'h80;
    mem[917] = 8'hff;
    mem[918] = 8'hff;
    mem[919] = 8'h03;
    mem[920] = 8'h00;
    mem[921] = 8'h00;
    mem[922] = 8'h00;
    mem[923] = 8'h00;
    mem[924] = 8'h00;
    mem[925] = 8'h00;
    mem[926] = 8'hf0;
    mem[927] = 8'h7f;
    mem[928] = 8'hfe;
    mem[929] = 8'h0f;
    mem[930] = 8'h00;
    mem[931] = 8'h00;
    mem[932] = 8'h80;
    mem[933] = 8'hff;
    mem[934] = 8'hff;
    mem[935] = 8'hff;
    mem[936] = 8'hff;
    mem[937] = 8'hff;
    mem[938] = 8'hff;
    mem[939] = 8'hff;
    mem[940] = 8'hff;
    mem[941] = 8'h01;
    mem[942] = 8'hf0;
    mem[943] = 8'h7f;
    mem[944] = 8'hfe;
    mem[945] = 8'h0f;
    mem[946] = 8'h00;
    mem[947] = 8'h00;
    mem[948] = 8'h80;
    mem[949] = 8'hff;
    mem[950] = 8'hff;
    mem[951] = 8'hff;
    mem[952] = 8'hff;
    mem[953] = 8'hff;
    mem[954] = 8'hff;
    mem[955] = 8'hff;
    mem[956] = 8'hff;
    mem[957] = 8'h01;
    mem[958] = 8'hf0;
    mem[959] = 8'h7f;
    mem[960] = 8'hfe;
    mem[961] = 8'h0f;
    mem[962] = 8'h00;
    mem[963] = 8'h00;
    mem[964] = 8'h80;
    mem[965] = 8'hff;
    mem[966] = 8'hff;
    mem[967] = 8'hff;
    mem[968] = 8'hff;
    mem[969] = 8'hff;
    mem[970] = 8'hff;
    mem[971] = 8'hff;
    mem[972] = 8'hff;
    mem[973] = 8'h01;
    mem[974] = 8'hf0;
    mem[975] = 8'h7f;
    mem[976] = 8'hfe;
    mem[977] = 8'h07;
    mem[978] = 8'h00;
    mem[979] = 8'h00;
    mem[980] = 8'h80;
    mem[981] = 8'hff;
    mem[982] = 8'hff;
    mem[983] = 8'hff;
    mem[984] = 8'hff;
    mem[985] = 8'hff;
    mem[986] = 8'hff;
    mem[987] = 8'hff;
    mem[988] = 8'hff;
    mem[989] = 8'h01;
    mem[990] = 8'hf0;
    mem[991] = 8'h7f;
    mem[992] = 8'hfe;
    mem[993] = 8'h07;
    mem[994] = 8'h00;
    mem[995] = 8'h00;
    mem[996] = 8'h80;
    mem[997] = 8'hff;
    mem[998] = 8'hff;
    mem[999] = 8'hff;
    mem[1000] = 8'hff;
    mem[1001] = 8'hff;
    mem[1002] = 8'hff;
    mem[1003] = 8'hff;
    mem[1004] = 8'hff;
    mem[1005] = 8'h01;
    mem[1006] = 8'hf0;
    mem[1007] = 8'h7f;
    mem[1008] = 8'hfe;
    mem[1009] = 8'h07;
    mem[1010] = 8'h00;
    mem[1011] = 8'h00;
    mem[1012] = 8'h80;
    mem[1013] = 8'hff;
    mem[1014] = 8'hff;
    mem[1015] = 8'hff;
    mem[1016] = 8'hff;
    mem[1017] = 8'hff;
    mem[1018] = 8'hff;
    mem[1019] = 8'hff;
    mem[1020] = 8'hff;
    mem[1021] = 8'h01;
    mem[1022] = 8'he0;
    mem[1023] = 8'h7f;
    mem[1024] = 8'hfe;
    mem[1025] = 8'h07;
    mem[1026] = 8'h00;
    mem[1027] = 8'h00;
    mem[1028] = 8'h80;
    mem[1029] = 8'hff;
    mem[1030] = 8'hff;
    mem[1031] = 8'hff;
    mem[1032] = 8'hff;
    mem[1033] = 8'hff;
    mem[1034] = 8'hff;
    mem[1035] = 8'hff;
    mem[1036] = 8'hff;
    mem[1037] = 8'h01;
    mem[1038] = 8'he0;
    mem[1039] = 8'h7f;
    mem[1040] = 8'hfe;
    mem[1041] = 8'h07;
    mem[1042] = 8'h00;
    mem[1043] = 8'h00;
    mem[1044] = 8'h80;
    mem[1045] = 8'hff;
    mem[1046] = 8'hff;
    mem[1047] = 8'hff;
    mem[1048] = 8'hff;
    mem[1049] = 8'hff;
    mem[1050] = 8'hff;
    mem[1051] = 8'hff;
    mem[1052] = 8'hff;
    mem[1053] = 8'h01;
    mem[1054] = 8'he0;
    mem[1055] = 8'h7f;
    mem[1056] = 8'hfe;
    mem[1057] = 8'h0f;
    mem[1058] = 8'h00;
    mem[1059] = 8'h00;
    mem[1060] = 8'h80;
    mem[1061] = 8'hff;
    mem[1062] = 8'hff;
    mem[1063] = 8'hff;
    mem[1064] = 8'hff;
    mem[1065] = 8'hff;
    mem[1066] = 8'hff;
    mem[1067] = 8'hff;
    mem[1068] = 8'hff;
    mem[1069] = 8'h01;
    mem[1070] = 8'hf0;
    mem[1071] = 8'h7f;
    mem[1072] = 8'hfe;
    mem[1073] = 8'h0f;
    mem[1074] = 8'h00;
    mem[1075] = 8'h00;
    mem[1076] = 8'h80;
    mem[1077] = 8'hff;
    mem[1078] = 8'hff;
    mem[1079] = 8'hff;
    mem[1080] = 8'hff;
    mem[1081] = 8'hff;
    mem[1082] = 8'hff;
    mem[1083] = 8'hff;
    mem[1084] = 8'hff;
    mem[1085] = 8'h01;
    mem[1086] = 8'hf0;
    mem[1087] = 8'h7f;
    mem[1088] = 8'hfe;
    mem[1089] = 8'h0f;
    mem[1090] = 8'h00;
    mem[1091] = 8'h00;
    mem[1092] = 8'h80;
    mem[1093] = 8'hff;
    mem[1094] = 8'hff;
    mem[1095] = 8'hff;
    mem[1096] = 8'hff;
    mem[1097] = 8'hff;
    mem[1098] = 8'hff;
    mem[1099] = 8'hff;
    mem[1100] = 8'hff;
    mem[1101] = 8'h01;
    mem[1102] = 8'hf0;
    mem[1103] = 8'h7f;
    mem[1104] = 8'hfe;
    mem[1105] = 8'h0f;
    mem[1106] = 8'h00;
    mem[1107] = 8'h00;
    mem[1108] = 8'h80;
    mem[1109] = 8'hff;
    mem[1110] = 8'hff;
    mem[1111] = 8'hff;
    mem[1112] = 8'hff;
    mem[1113] = 8'hff;
    mem[1114] = 8'hff;
    mem[1115] = 8'hff;
    mem[1116] = 8'hff;
    mem[1117] = 8'h01;
    mem[1118] = 8'hf0;
    mem[1119] = 8'h7f;
    mem[1120] = 8'hfe;
    mem[1121] = 8'h0f;
    mem[1122] = 8'h00;
    mem[1123] = 8'h00;
    mem[1124] = 8'h80;
    mem[1125] = 8'hff;
    mem[1126] = 8'hff;
    mem[1127] = 8'hff;
    mem[1128] = 8'hff;
    mem[1129] = 8'hff;
    mem[1130] = 8'hff;
    mem[1131] = 8'hff;
    mem[1132] = 8'hff;
    mem[1133] = 8'h01;
    mem[1134] = 8'hf0;
    mem[1135] = 8'h7f;
    mem[1136] = 8'hfe;
    mem[1137] = 8'h0f;
    mem[1138] = 8'h00;
    mem[1139] = 8'h00;
    mem[1140] = 8'h80;
    mem[1141] = 8'hff;
    mem[1142] = 8'hff;
    mem[1143] = 8'hff;
    mem[1144] = 8'hff;
    mem[1145] = 8'hff;
    mem[1146] = 8'hff;
    mem[1147] = 8'hff;
    mem[1148] = 8'hff;
    mem[1149] = 8'h01;
    mem[1150] = 8'hf0;
    mem[1151] = 8'h7f;
    mem[1152] = 8'hfe;
    mem[1153] = 8'h0f;
    mem[1154] = 8'h00;
    mem[1155] = 8'h00;
    mem[1156] = 8'h80;
    mem[1157] = 8'hff;
    mem[1158] = 8'hff;
    mem[1159] = 8'hff;
    mem[1160] = 8'hff;
    mem[1161] = 8'hff;
    mem[1162] = 8'hff;
    mem[1163] = 8'hff;
    mem[1164] = 8'hff;
    mem[1165] = 8'h01;
    mem[1166] = 8'hf0;
    mem[1167] = 8'h7f;
    mem[1168] = 8'hfc;
    mem[1169] = 8'h0f;
    mem[1170] = 8'h00;
    mem[1171] = 8'h00;
    mem[1172] = 8'h80;
    mem[1173] = 8'hff;
    mem[1174] = 8'hff;
    mem[1175] = 8'hff;
    mem[1176] = 8'hff;
    mem[1177] = 8'hff;
    mem[1178] = 8'hff;
    mem[1179] = 8'hff;
    mem[1180] = 8'hff;
    mem[1181] = 8'h01;
    mem[1182] = 8'hf0;
    mem[1183] = 8'h3f;
    mem[1184] = 8'hfc;
    mem[1185] = 8'h1f;
    mem[1186] = 8'h00;
    mem[1187] = 8'h00;
    mem[1188] = 8'h80;
    mem[1189] = 8'hff;
    mem[1190] = 8'hff;
    mem[1191] = 8'hff;
    mem[1192] = 8'hff;
    mem[1193] = 8'hff;
    mem[1194] = 8'hff;
    mem[1195] = 8'hff;
    mem[1196] = 8'hff;
    mem[1197] = 8'h01;
    mem[1198] = 8'hf8;
    mem[1199] = 8'h3f;
    mem[1200] = 8'hfc;
    mem[1201] = 8'h1f;
    mem[1202] = 8'h00;
    mem[1203] = 8'h00;
    mem[1204] = 8'h80;
    mem[1205] = 8'hff;
    mem[1206] = 8'hff;
    mem[1207] = 8'hff;
    mem[1208] = 8'hff;
    mem[1209] = 8'hff;
    mem[1210] = 8'hff;
    mem[1211] = 8'hff;
    mem[1212] = 8'hff;
    mem[1213] = 8'h01;
    mem[1214] = 8'hf8;
    mem[1215] = 8'h3f;
    mem[1216] = 8'hfc;
    mem[1217] = 8'h1f;
    mem[1218] = 8'h00;
    mem[1219] = 8'h00;
    mem[1220] = 8'h80;
    mem[1221] = 8'hff;
    mem[1222] = 8'hff;
    mem[1223] = 8'h03;
    mem[1224] = 8'hf0;
    mem[1225] = 8'hff;
    mem[1226] = 8'h7f;
    mem[1227] = 8'h00;
    mem[1228] = 8'h00;
    mem[1229] = 8'h00;
    mem[1230] = 8'hf8;
    mem[1231] = 8'h3f;
    mem[1232] = 8'hfc;
    mem[1233] = 8'h1f;
    mem[1234] = 8'h00;
    mem[1235] = 8'h00;
    mem[1236] = 8'h80;
    mem[1237] = 8'hff;
    mem[1238] = 8'hff;
    mem[1239] = 8'h03;
    mem[1240] = 8'hf0;
    mem[1241] = 8'hff;
    mem[1242] = 8'h7f;
    mem[1243] = 8'h00;
    mem[1244] = 8'h00;
    mem[1245] = 8'h00;
    mem[1246] = 8'hf8;
    mem[1247] = 8'h3f;
    mem[1248] = 8'hfc;
    mem[1249] = 8'h3f;
    mem[1250] = 8'h00;
    mem[1251] = 8'h00;
    mem[1252] = 8'h80;
    mem[1253] = 8'hff;
    mem[1254] = 8'hff;
    mem[1255] = 8'h03;
    mem[1256] = 8'hf0;
    mem[1257] = 8'hff;
    mem[1258] = 8'h7f;
    mem[1259] = 8'h00;
    mem[1260] = 8'h00;
    mem[1261] = 8'h00;
    mem[1262] = 8'hfc;
    mem[1263] = 8'h3f;
    mem[1264] = 8'hf8;
    mem[1265] = 8'h3f;
    mem[1266] = 8'h00;
    mem[1267] = 8'h00;
    mem[1268] = 8'h80;
    mem[1269] = 8'hff;
    mem[1270] = 8'hff;
    mem[1271] = 8'h03;
    mem[1272] = 8'hf0;
    mem[1273] = 8'hff;
    mem[1274] = 8'h7f;
    mem[1275] = 8'h00;
    mem[1276] = 8'h00;
    mem[1277] = 8'h00;
    mem[1278] = 8'hfc;
    mem[1279] = 8'h1f;
    mem[1280] = 8'hf8;
    mem[1281] = 8'h3f;
    mem[1282] = 8'h00;
    mem[1283] = 8'h00;
    mem[1284] = 8'h80;
    mem[1285] = 8'hff;
    mem[1286] = 8'hff;
    mem[1287] = 8'h03;
    mem[1288] = 8'hf0;
    mem[1289] = 8'hff;
    mem[1290] = 8'h7f;
    mem[1291] = 8'h00;
    mem[1292] = 8'h00;
    mem[1293] = 8'h00;
    mem[1294] = 8'hfc;
    mem[1295] = 8'h1f;
    mem[1296] = 8'hf8;
    mem[1297] = 8'h7f;
    mem[1298] = 8'h00;
    mem[1299] = 8'h00;
    mem[1300] = 8'h80;
    mem[1301] = 8'hff;
    mem[1302] = 8'hff;
    mem[1303] = 8'h03;
    mem[1304] = 8'hf0;
    mem[1305] = 8'hff;
    mem[1306] = 8'h7f;
    mem[1307] = 8'h00;
    mem[1308] = 8'h00;
    mem[1309] = 8'h00;
    mem[1310] = 8'hfe;
    mem[1311] = 8'h1f;
    mem[1312] = 8'hf0;
    mem[1313] = 8'h7f;
    mem[1314] = 8'h00;
    mem[1315] = 8'h00;
    mem[1316] = 8'h80;
    mem[1317] = 8'hff;
    mem[1318] = 8'hff;
    mem[1319] = 8'h03;
    mem[1320] = 8'hf0;
    mem[1321] = 8'hff;
    mem[1322] = 8'h7f;
    mem[1323] = 8'h00;
    mem[1324] = 8'h00;
    mem[1325] = 8'h00;
    mem[1326] = 8'hfe;
    mem[1327] = 8'h0f;
    mem[1328] = 8'hf0;
    mem[1329] = 8'h7f;
    mem[1330] = 8'h00;
    mem[1331] = 8'h00;
    mem[1332] = 8'h80;
    mem[1333] = 8'hff;
    mem[1334] = 8'hff;
    mem[1335] = 8'h03;
    mem[1336] = 8'hf0;
    mem[1337] = 8'hff;
    mem[1338] = 8'h7f;
    mem[1339] = 8'h00;
    mem[1340] = 8'h00;
    mem[1341] = 8'h00;
    mem[1342] = 8'hfe;
    mem[1343] = 8'h0f;
    mem[1344] = 8'hf0;
    mem[1345] = 8'hff;
    mem[1346] = 8'h00;
    mem[1347] = 8'h00;
    mem[1348] = 8'h80;
    mem[1349] = 8'hff;
    mem[1350] = 8'hff;
    mem[1351] = 8'h03;
    mem[1352] = 8'hf0;
    mem[1353] = 8'hff;
    mem[1354] = 8'h7f;
    mem[1355] = 8'h00;
    mem[1356] = 8'h00;
    mem[1357] = 8'h00;
    mem[1358] = 8'hff;
    mem[1359] = 8'h0f;
    mem[1360] = 8'he0;
    mem[1361] = 8'hff;
    mem[1362] = 8'h00;
    mem[1363] = 8'h00;
    mem[1364] = 8'h80;
    mem[1365] = 8'hff;
    mem[1366] = 8'hff;
    mem[1367] = 8'h03;
    mem[1368] = 8'hf0;
    mem[1369] = 8'hff;
    mem[1370] = 8'h7f;
    mem[1371] = 8'h00;
    mem[1372] = 8'h00;
    mem[1373] = 8'h00;
    mem[1374] = 8'hff;
    mem[1375] = 8'h07;
    mem[1376] = 8'he0;
    mem[1377] = 8'hff;
    mem[1378] = 8'h01;
    mem[1379] = 8'h00;
    mem[1380] = 8'h80;
    mem[1381] = 8'hff;
    mem[1382] = 8'hff;
    mem[1383] = 8'h03;
    mem[1384] = 8'hf0;
    mem[1385] = 8'hff;
    mem[1386] = 8'h7f;
    mem[1387] = 8'h00;
    mem[1388] = 8'h00;
    mem[1389] = 8'h80;
    mem[1390] = 8'hff;
    mem[1391] = 8'h07;
    mem[1392] = 8'he0;
    mem[1393] = 8'hff;
    mem[1394] = 8'h01;
    mem[1395] = 8'h00;
    mem[1396] = 8'h00;
    mem[1397] = 8'h00;
    mem[1398] = 8'h00;
    mem[1399] = 8'h00;
    mem[1400] = 8'hf0;
    mem[1401] = 8'hff;
    mem[1402] = 8'h7f;
    mem[1403] = 8'h00;
    mem[1404] = 8'h00;
    mem[1405] = 8'h80;
    mem[1406] = 8'hff;
    mem[1407] = 8'h07;
    mem[1408] = 8'hc0;
    mem[1409] = 8'hff;
    mem[1410] = 8'h03;
    mem[1411] = 8'h00;
    mem[1412] = 8'h00;
    mem[1413] = 8'h00;
    mem[1414] = 8'h00;
    mem[1415] = 8'h00;
    mem[1416] = 8'hf0;
    mem[1417] = 8'hff;
    mem[1418] = 8'h7f;
    mem[1419] = 8'h00;
    mem[1420] = 8'h00;
    mem[1421] = 8'hc0;
    mem[1422] = 8'hff;
    mem[1423] = 8'h03;
    mem[1424] = 8'hc0;
    mem[1425] = 8'hff;
    mem[1426] = 8'h03;
    mem[1427] = 8'h00;
    mem[1428] = 8'h00;
    mem[1429] = 8'h00;
    mem[1430] = 8'h00;
    mem[1431] = 8'h00;
    mem[1432] = 8'hf0;
    mem[1433] = 8'hff;
    mem[1434] = 8'h7f;
    mem[1435] = 8'h00;
    mem[1436] = 8'h00;
    mem[1437] = 8'hc0;
    mem[1438] = 8'hff;
    mem[1439] = 8'h03;
    mem[1440] = 8'h80;
    mem[1441] = 8'hff;
    mem[1442] = 8'h07;
    mem[1443] = 8'h00;
    mem[1444] = 8'h00;
    mem[1445] = 8'h00;
    mem[1446] = 8'h00;
    mem[1447] = 8'h00;
    mem[1448] = 8'hf0;
    mem[1449] = 8'hff;
    mem[1450] = 8'h7f;
    mem[1451] = 8'h00;
    mem[1452] = 8'h00;
    mem[1453] = 8'he0;
    mem[1454] = 8'hff;
    mem[1455] = 8'h01;
    mem[1456] = 8'h80;
    mem[1457] = 8'hff;
    mem[1458] = 8'h07;
    mem[1459] = 8'h00;
    mem[1460] = 8'h00;
    mem[1461] = 8'h00;
    mem[1462] = 8'h00;
    mem[1463] = 8'h00;
    mem[1464] = 8'hf0;
    mem[1465] = 8'hff;
    mem[1466] = 8'h7f;
    mem[1467] = 8'h00;
    mem[1468] = 8'h00;
    mem[1469] = 8'he0;
    mem[1470] = 8'hff;
    mem[1471] = 8'h01;
    mem[1472] = 8'h00;
    mem[1473] = 8'hff;
    mem[1474] = 8'h0f;
    mem[1475] = 8'h00;
    mem[1476] = 8'h00;
    mem[1477] = 8'h00;
    mem[1478] = 8'h00;
    mem[1479] = 8'h00;
    mem[1480] = 8'hf0;
    mem[1481] = 8'hff;
    mem[1482] = 8'h7f;
    mem[1483] = 8'h00;
    mem[1484] = 8'h00;
    mem[1485] = 8'hf0;
    mem[1486] = 8'hff;
    mem[1487] = 8'h00;
    mem[1488] = 8'h00;
    mem[1489] = 8'hff;
    mem[1490] = 8'h1f;
    mem[1491] = 8'h00;
    mem[1492] = 8'h00;
    mem[1493] = 8'h00;
    mem[1494] = 8'h00;
    mem[1495] = 8'h00;
    mem[1496] = 8'hf0;
    mem[1497] = 8'hff;
    mem[1498] = 8'h7f;
    mem[1499] = 8'h00;
    mem[1500] = 8'h00;
    mem[1501] = 8'hf8;
    mem[1502] = 8'hff;
    mem[1503] = 8'h00;
    mem[1504] = 8'h00;
    mem[1505] = 8'hfe;
    mem[1506] = 8'h1f;
    mem[1507] = 8'h00;
    mem[1508] = 8'h00;
    mem[1509] = 8'h00;
    mem[1510] = 8'h00;
    mem[1511] = 8'h00;
    mem[1512] = 8'hf0;
    mem[1513] = 8'hff;
    mem[1514] = 8'h7f;
    mem[1515] = 8'h00;
    mem[1516] = 8'h00;
    mem[1517] = 8'hf8;
    mem[1518] = 8'h7f;
    mem[1519] = 8'h00;
    mem[1520] = 8'h00;
    mem[1521] = 8'hfe;
    mem[1522] = 8'h3f;
    mem[1523] = 8'h00;
    mem[1524] = 8'h00;
    mem[1525] = 8'h00;
    mem[1526] = 8'h00;
    mem[1527] = 8'h00;
    mem[1528] = 8'hf0;
    mem[1529] = 8'hff;
    mem[1530] = 8'h7f;
    mem[1531] = 8'h00;
    mem[1532] = 8'h00;
    mem[1533] = 8'hfc;
    mem[1534] = 8'h7f;
    mem[1535] = 8'h00;
    mem[1536] = 8'h00;
    mem[1537] = 8'hfc;
    mem[1538] = 8'h7f;
    mem[1539] = 8'h00;
    mem[1540] = 8'h00;
    mem[1541] = 8'h00;
    mem[1542] = 8'h00;
    mem[1543] = 8'h00;
    mem[1544] = 8'hf0;
    mem[1545] = 8'hff;
    mem[1546] = 8'h7f;
    mem[1547] = 8'h00;
    mem[1548] = 8'h00;
    mem[1549] = 8'hfe;
    mem[1550] = 8'h3f;
    mem[1551] = 8'h00;
    mem[1552] = 8'h00;
    mem[1553] = 8'hfc;
    mem[1554] = 8'hff;
    mem[1555] = 8'h00;
    mem[1556] = 8'h00;
    mem[1557] = 8'h00;
    mem[1558] = 8'h00;
    mem[1559] = 8'h00;
    mem[1560] = 8'hf0;
    mem[1561] = 8'hff;
    mem[1562] = 8'h7f;
    mem[1563] = 8'h00;
    mem[1564] = 8'h00;
    mem[1565] = 8'hff;
    mem[1566] = 8'h3f;
    mem[1567] = 8'h00;
    mem[1568] = 8'h00;
    mem[1569] = 8'hf8;
    mem[1570] = 8'hff;
    mem[1571] = 8'h01;
    mem[1572] = 8'h00;
    mem[1573] = 8'h00;
    mem[1574] = 8'h00;
    mem[1575] = 8'h00;
    mem[1576] = 8'hf0;
    mem[1577] = 8'hff;
    mem[1578] = 8'h7f;
    mem[1579] = 8'h00;
    mem[1580] = 8'h80;
    mem[1581] = 8'hff;
    mem[1582] = 8'h1f;
    mem[1583] = 8'h00;
    mem[1584] = 8'h00;
    mem[1585] = 8'hf0;
    mem[1586] = 8'hff;
    mem[1587] = 8'h03;
    mem[1588] = 8'h00;
    mem[1589] = 8'h00;
    mem[1590] = 8'h00;
    mem[1591] = 8'h00;
    mem[1592] = 8'hf0;
    mem[1593] = 8'hff;
    mem[1594] = 8'h7f;
    mem[1595] = 8'h00;
    mem[1596] = 8'hc0;
    mem[1597] = 8'hff;
    mem[1598] = 8'h0f;
    mem[1599] = 8'h00;
    mem[1600] = 8'h00;
    mem[1601] = 8'hf0;
    mem[1602] = 8'hff;
    mem[1603] = 8'h03;
    mem[1604] = 8'h00;
    mem[1605] = 8'h00;
    mem[1606] = 8'h00;
    mem[1607] = 8'h00;
    mem[1608] = 8'hf0;
    mem[1609] = 8'hff;
    mem[1610] = 8'h7f;
    mem[1611] = 8'h00;
    mem[1612] = 8'hc0;
    mem[1613] = 8'hff;
    mem[1614] = 8'h0f;
    mem[1615] = 8'h00;
    mem[1616] = 8'h00;
    mem[1617] = 8'he0;
    mem[1618] = 8'hff;
    mem[1619] = 8'h07;
    mem[1620] = 8'h00;
    mem[1621] = 8'h00;
    mem[1622] = 8'h00;
    mem[1623] = 8'h00;
    mem[1624] = 8'hf0;
    mem[1625] = 8'hff;
    mem[1626] = 8'h7f;
    mem[1627] = 8'h00;
    mem[1628] = 8'he0;
    mem[1629] = 8'hff;
    mem[1630] = 8'h07;
    mem[1631] = 8'h00;
    mem[1632] = 8'h00;
    mem[1633] = 8'hc0;
    mem[1634] = 8'hff;
    mem[1635] = 8'h1f;
    mem[1636] = 8'h00;
    mem[1637] = 8'h00;
    mem[1638] = 8'h00;
    mem[1639] = 8'h00;
    mem[1640] = 8'hf0;
    mem[1641] = 8'hff;
    mem[1642] = 8'h7f;
    mem[1643] = 8'h00;
    mem[1644] = 8'hf0;
    mem[1645] = 8'hff;
    mem[1646] = 8'h03;
    mem[1647] = 8'h00;
    mem[1648] = 8'h00;
    mem[1649] = 8'h80;
    mem[1650] = 8'hff;
    mem[1651] = 8'h3f;
    mem[1652] = 8'h00;
    mem[1653] = 8'h00;
    mem[1654] = 8'h00;
    mem[1655] = 8'h00;
    mem[1656] = 8'hf0;
    mem[1657] = 8'hff;
    mem[1658] = 8'h7f;
    mem[1659] = 8'h00;
    mem[1660] = 8'hfc;
    mem[1661] = 8'hff;
    mem[1662] = 8'h01;
    mem[1663] = 8'h00;
    mem[1664] = 8'h00;
    mem[1665] = 8'h80;
    mem[1666] = 8'hff;
    mem[1667] = 8'h7f;
    mem[1668] = 8'h00;
    mem[1669] = 8'h00;
    mem[1670] = 8'h00;
    mem[1671] = 8'h00;
    mem[1672] = 8'hf0;
    mem[1673] = 8'hff;
    mem[1674] = 8'h7f;
    mem[1675] = 8'h00;
    mem[1676] = 8'hfe;
    mem[1677] = 8'hff;
    mem[1678] = 8'h01;
    mem[1679] = 8'h00;
    mem[1680] = 8'h00;
    mem[1681] = 8'h00;
    mem[1682] = 8'hff;
    mem[1683] = 8'hff;
    mem[1684] = 8'h00;
    mem[1685] = 8'h00;
    mem[1686] = 8'h00;
    mem[1687] = 8'h00;
    mem[1688] = 8'hf0;
    mem[1689] = 8'hff;
    mem[1690] = 8'h7f;
    mem[1691] = 8'h00;
    mem[1692] = 8'hff;
    mem[1693] = 8'hff;
    mem[1694] = 8'h00;
    mem[1695] = 8'h00;
    mem[1696] = 8'h00;
    mem[1697] = 8'h00;
    mem[1698] = 8'hfe;
    mem[1699] = 8'hff;
    mem[1700] = 8'h01;
    mem[1701] = 8'h00;
    mem[1702] = 8'h00;
    mem[1703] = 8'h00;
    mem[1704] = 8'hf0;
    mem[1705] = 8'hff;
    mem[1706] = 8'h7f;
    mem[1707] = 8'h80;
    mem[1708] = 8'hff;
    mem[1709] = 8'h7f;
    mem[1710] = 8'h00;
    mem[1711] = 8'h00;
    mem[1712] = 8'h00;
    mem[1713] = 8'h00;
    mem[1714] = 8'hfc;
    mem[1715] = 8'hff;
    mem[1716] = 8'h07;
    mem[1717] = 8'h00;
    mem[1718] = 8'h00;
    mem[1719] = 8'h00;
    mem[1720] = 8'hf0;
    mem[1721] = 8'hff;
    mem[1722] = 8'h7f;
    mem[1723] = 8'he0;
    mem[1724] = 8'hff;
    mem[1725] = 8'h3f;
    mem[1726] = 8'h00;
    mem[1727] = 8'h00;
    mem[1728] = 8'h00;
    mem[1729] = 8'h00;
    mem[1730] = 8'hf8;
    mem[1731] = 8'hff;
    mem[1732] = 8'h0f;
    mem[1733] = 8'h00;
    mem[1734] = 8'h00;
    mem[1735] = 8'h00;
    mem[1736] = 8'hf0;
    mem[1737] = 8'hff;
    mem[1738] = 8'h7f;
    mem[1739] = 8'hf0;
    mem[1740] = 8'hff;
    mem[1741] = 8'h1f;
    mem[1742] = 8'h00;
    mem[1743] = 8'h00;
    mem[1744] = 8'h00;
    mem[1745] = 8'h00;
    mem[1746] = 8'hf0;
    mem[1747] = 8'hff;
    mem[1748] = 8'h3f;
    mem[1749] = 8'h00;
    mem[1750] = 8'h00;
    mem[1751] = 8'h00;
    mem[1752] = 8'hf0;
    mem[1753] = 8'hff;
    mem[1754] = 8'h7f;
    mem[1755] = 8'hf0;
    mem[1756] = 8'hff;
    mem[1757] = 8'h0f;
    mem[1758] = 8'h00;
    mem[1759] = 8'h00;
    mem[1760] = 8'h00;
    mem[1761] = 8'h00;
    mem[1762] = 8'he0;
    mem[1763] = 8'hff;
    mem[1764] = 8'hff;
    mem[1765] = 8'h00;
    mem[1766] = 8'h00;
    mem[1767] = 8'h00;
    mem[1768] = 8'hf0;
    mem[1769] = 8'hff;
    mem[1770] = 8'h7f;
    mem[1771] = 8'hf0;
    mem[1772] = 8'hff;
    mem[1773] = 8'h07;
    mem[1774] = 8'h00;
    mem[1775] = 8'h00;
    mem[1776] = 8'h00;
    mem[1777] = 8'h00;
    mem[1778] = 8'hc0;
    mem[1779] = 8'hff;
    mem[1780] = 8'hff;
    mem[1781] = 8'h03;
    mem[1782] = 8'h00;
    mem[1783] = 8'h00;
    mem[1784] = 8'hf0;
    mem[1785] = 8'hff;
    mem[1786] = 8'h7f;
    mem[1787] = 8'hf0;
    mem[1788] = 8'hff;
    mem[1789] = 8'h03;
    mem[1790] = 8'h00;
    mem[1791] = 8'h00;
    mem[1792] = 8'h00;
    mem[1793] = 8'h00;
    mem[1794] = 8'h80;
    mem[1795] = 8'hff;
    mem[1796] = 8'hff;
    mem[1797] = 8'h0f;
    mem[1798] = 8'h00;
    mem[1799] = 8'h00;
    mem[1800] = 8'hf0;
    mem[1801] = 8'hff;
    mem[1802] = 8'h7f;
    mem[1803] = 8'hf0;
    mem[1804] = 8'hff;
    mem[1805] = 8'h01;
    mem[1806] = 8'h00;
    mem[1807] = 8'h00;
    mem[1808] = 8'h00;
    mem[1809] = 8'h00;
    mem[1810] = 8'h00;
    mem[1811] = 8'hfe;
    mem[1812] = 8'hff;
    mem[1813] = 8'h7f;
    mem[1814] = 8'h00;
    mem[1815] = 8'h00;
    mem[1816] = 8'hf0;
    mem[1817] = 8'hff;
    mem[1818] = 8'h7f;
    mem[1819] = 8'hf0;
    mem[1820] = 8'h7f;
    mem[1821] = 8'h00;
    mem[1822] = 8'h00;
    mem[1823] = 8'h00;
    mem[1824] = 8'h00;
    mem[1825] = 8'h00;
    mem[1826] = 8'h00;
    mem[1827] = 8'hfc;
    mem[1828] = 8'hff;
    mem[1829] = 8'hff;
    mem[1830] = 8'h03;
    mem[1831] = 8'h00;
    mem[1832] = 8'hf0;
    mem[1833] = 8'hff;
    mem[1834] = 8'h7f;
    mem[1835] = 8'hf0;
    mem[1836] = 8'h3f;
    mem[1837] = 8'h00;
    mem[1838] = 8'h00;
    mem[1839] = 8'h00;
    mem[1840] = 8'h00;
    mem[1841] = 8'h00;
    mem[1842] = 8'h00;
    mem[1843] = 8'hf8;
    mem[1844] = 8'hff;
    mem[1845] = 8'hff;
    mem[1846] = 8'h3f;
    mem[1847] = 8'h00;
    mem[1848] = 8'hf0;
    mem[1849] = 8'hff;
    mem[1850] = 8'h7f;
    mem[1851] = 8'hf0;
    mem[1852] = 8'h1f;
    mem[1853] = 8'h00;
    mem[1854] = 8'h00;
    mem[1855] = 8'h00;
    mem[1856] = 8'h00;
    mem[1857] = 8'h00;
    mem[1858] = 8'h00;
    mem[1859] = 8'he0;
    mem[1860] = 8'hff;
    mem[1861] = 8'hff;
    mem[1862] = 8'hff;
    mem[1863] = 8'h7f;
    mem[1864] = 8'hfc;
    mem[1865] = 8'hff;
    mem[1866] = 8'h7f;
    mem[1867] = 8'hf0;
    mem[1868] = 8'h07;
    mem[1869] = 8'h00;
    mem[1870] = 8'h00;
    mem[1871] = 8'h00;
    mem[1872] = 8'h00;
    mem[1873] = 8'h00;
    mem[1874] = 8'h00;
    mem[1875] = 8'hc0;
    mem[1876] = 8'hff;
    mem[1877] = 8'hff;
    mem[1878] = 8'hff;
    mem[1879] = 8'hff;
    mem[1880] = 8'hff;
    mem[1881] = 8'hff;
    mem[1882] = 8'h7f;
    mem[1883] = 8'hf0;
    mem[1884] = 8'h03;
    mem[1885] = 8'h00;
    mem[1886] = 8'h00;
    mem[1887] = 8'h00;
    mem[1888] = 8'h00;
    mem[1889] = 8'h00;
    mem[1890] = 8'h00;
    mem[1891] = 8'h00;
    mem[1892] = 8'hff;
    mem[1893] = 8'hff;
    mem[1894] = 8'hff;
    mem[1895] = 8'hff;
    mem[1896] = 8'hff;
    mem[1897] = 8'hff;
    mem[1898] = 8'h7f;
    mem[1899] = 8'hf0;
    mem[1900] = 8'h00;
    mem[1901] = 8'h00;
    mem[1902] = 8'h00;
    mem[1903] = 8'h00;
    mem[1904] = 8'h00;
    mem[1905] = 8'h00;
    mem[1906] = 8'h00;
    mem[1907] = 8'h00;
    mem[1908] = 8'hfc;
    mem[1909] = 8'hff;
    mem[1910] = 8'hff;
    mem[1911] = 8'hff;
    mem[1912] = 8'hff;
    mem[1913] = 8'hff;
    mem[1914] = 8'h7f;
    mem[1915] = 8'h30;
    mem[1916] = 8'h00;
    mem[1917] = 8'h00;
    mem[1918] = 8'h00;
    mem[1919] = 8'h00;
    mem[1920] = 8'h00;
    mem[1921] = 8'h00;
    mem[1922] = 8'h00;
    mem[1923] = 8'h00;
    mem[1924] = 8'hf0;
    mem[1925] = 8'hff;
    mem[1926] = 8'hff;
    mem[1927] = 8'hff;
    mem[1928] = 8'hff;
    mem[1929] = 8'hff;
    mem[1930] = 8'h7f;
    mem[1931] = 8'h00;
    mem[1932] = 8'h00;
    mem[1933] = 8'h00;
    mem[1934] = 8'h00;
    mem[1935] = 8'h00;
    mem[1936] = 8'h00;
    mem[1937] = 8'h00;
    mem[1938] = 8'h00;
    mem[1939] = 8'h00;
    mem[1940] = 8'hc0;
    mem[1941] = 8'hff;
    mem[1942] = 8'hff;
    mem[1943] = 8'hff;
    mem[1944] = 8'hff;
    mem[1945] = 8'hff;
    mem[1946] = 8'h7f;
    mem[1947] = 8'h00;
    mem[1948] = 8'h00;
    mem[1949] = 8'h00;
    mem[1950] = 8'h00;
    mem[1951] = 8'h00;
    mem[1952] = 8'h00;
    mem[1953] = 8'h00;
    mem[1954] = 8'h00;
    mem[1955] = 8'h00;
    mem[1956] = 8'h00;
    mem[1957] = 8'hff;
    mem[1958] = 8'hff;
    mem[1959] = 8'hff;
    mem[1960] = 8'hff;
    mem[1961] = 8'hff;
    mem[1962] = 8'h7f;
    mem[1963] = 8'h00;
    mem[1964] = 8'h00;
    mem[1965] = 8'h00;
    mem[1966] = 8'h00;
    mem[1967] = 8'h00;
    mem[1968] = 8'h00;
    mem[1969] = 8'h00;
    mem[1970] = 8'h00;
    mem[1971] = 8'h00;
    mem[1972] = 8'h00;
    mem[1973] = 8'hf8;
    mem[1974] = 8'hff;
    mem[1975] = 8'hff;
    mem[1976] = 8'hff;
    mem[1977] = 8'hff;
    mem[1978] = 8'h1f;
    mem[1979] = 8'h00;
    mem[1980] = 8'h00;
    mem[1981] = 8'h00;
    mem[1982] = 8'h00;
    mem[1983] = 8'h00;
    mem[1984] = 8'h00;
    mem[1985] = 8'h00;
    mem[1986] = 8'h00;
    mem[1987] = 8'h00;
    mem[1988] = 8'h00;
    mem[1989] = 8'hc0;
    mem[1990] = 8'hff;
    mem[1991] = 8'hff;
    mem[1992] = 8'hff;
    mem[1993] = 8'hff;
    mem[1994] = 8'h03;
    mem[1995] = 8'h00;
    mem[1996] = 8'h00;
    mem[1997] = 8'h00;
    mem[1998] = 8'h00;
    mem[1999] = 8'h00;
    mem[2000] = 8'h00;
    mem[2001] = 8'h00;
    mem[2002] = 8'h00;
    mem[2003] = 8'h00;
    mem[2004] = 8'h00;
    mem[2005] = 8'h00;
    mem[2006] = 8'hfc;
    mem[2007] = 8'hff;
    mem[2008] = 8'hff;
    mem[2009] = 8'h3f;
    mem[2010] = 8'h00;
    mem[2011] = 8'h00;
    mem[2012] = 8'h00;
    mem[2013] = 8'h00;
    mem[2014] = 8'h00;
    mem[2015] = 8'h00;
    mem[2016] = 8'h00;
    mem[2017] = 8'h00;
    mem[2018] = 8'h00;
    mem[2019] = 8'h00;
    mem[2020] = 8'h00;
    mem[2021] = 8'h00;
    mem[2022] = 8'h80;
    mem[2023] = 8'hff;
    mem[2024] = 8'hff;
    mem[2025] = 8'h01;
    mem[2026] = 8'h00;
    mem[2027] = 8'h00;
    mem[2028] = 8'h00;
    mem[2029] = 8'h00;
    mem[2030] = 8'h00;
    mem[2031] = 8'h00;
    mem[2032] = 8'h00;
    mem[2033] = 8'h00;
    mem[2034] = 8'h00;
    mem[2035] = 8'h00;
    mem[2036] = 8'h00;
    mem[2037] = 8'h00;
    mem[2038] = 8'h00;
    mem[2039] = 8'h00;
    mem[2040] = 8'h00;
    mem[2041] = 8'h00;
    mem[2042] = 8'h00;
    mem[2043] = 8'h00;
    mem[2044] = 8'h00;
    mem[2045] = 8'h00;
    mem[2046] = 8'h00;
    mem[2047] = 8'h00;
  end

  wire [10:0] addr = {y[6:0], x[6:3]};
  assign pixel = mem[addr][x&7];

endmodule
