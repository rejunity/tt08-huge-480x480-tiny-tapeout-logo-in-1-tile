/*
 * Copyright (c) 2024 Tiny Tapeout LTD
 * SPDX-License-Identifier: Apache-2.0
 * Author: Renaldas Zioma
 */

`default_nettype none

parameter LOGO_SIZE = 272;  // Size of the logo in pixels
parameter DISPLAY_WIDTH = 640;  // VGA display width
parameter DISPLAY_HEIGHT = 480;  // VGA display height

`define COLOR_WHITE 3'd7

module tt_um_rejunity_vga_logo (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // VGA signals
  wire hsync;
  wire vsync;
  reg [1:0] R;
  reg [1:0] G;
  reg [1:0] B;
  wire video_active;
  wire [9:0] pix_x;
  wire [9:0] pix_y;


  // TinyVGA PMOD
  assign uo_out  = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

  // Unused outputs assigned to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in[7:1], uio_in};

  hvsync_generator vga_sync_gen (
      .clk(clk),
      .reset(~rst_n),
      .hsync(hsync),
      .vsync(vsync),
      .display_on(video_active),
      .hpos(pix_x),
      .vpos(pix_y)
  );

  reg pixel_value;

  // bitmap_rom rom1 (
  //     .x(pix_x[6:0]),
  //     .y(pix_y[6:0]),
  //     .pixel(pixel_value)
  // );

  reg [11:0] addr;
  reg [7:0] len;
  bitmap_rom_rle rom2 (
    .addr(addr),
    .len(len)
  );

  assign {R, G, B } = video_active*pixel_value*6'b11_11_00;

  // increase couner every frame (vsync happens once per frame)
  reg [11:0] counter;
  always @(posedge clk) begin
    if (~rst_n) begin
      counter <= 0;
    end else begin
      if (vsync) begin
        addr <= 0;
        counter <= 0;
        pixel_value <= 0;
      end else if (pix_x < LOGO_SIZE && pix_y < LOGO_SIZE) begin
        if (counter >= len) begin
          addr <= addr + 1;
          counter <= 0;
          pixel_value <= ~pixel_value;
        end else
          counter <= counter + 1;
      end
    end
  end  

endmodule

// --------------------------------------------------------

module bitmap_rom_rle (
    input wire [11:0] addr,
    output wire [7:0] len
);

  reg [7:0] mem[1329:0];
  initial begin
    mem[11'h000] = 8'h87;
    mem[11'h001] = 8'h01;
    mem[11'h002] = 8'hfd;
    mem[11'h003] = 8'h21;
    mem[11'h004] = 8'he7;
    mem[11'h005] = 8'h2d;
    mem[11'h006] = 8'hdc;
    mem[11'h007] = 8'h38;
    mem[11'h008] = 8'hd1;
    mem[11'h009] = 8'h41;
    mem[11'h00a] = 8'hca;
    mem[11'h00b] = 8'h48;
    mem[11'h00c] = 8'hc2;
    mem[11'h00d] = 8'h4f;
    mem[11'h00e] = 8'hbc;
    mem[11'h00f] = 8'h55;
    mem[11'h010] = 8'hb6;
    mem[11'h011] = 8'h5b;
    mem[11'h012] = 8'hb0;
    mem[11'h013] = 8'h61;
    mem[11'h014] = 8'hab;
    mem[11'h015] = 8'h65;
    mem[11'h016] = 8'ha7;
    mem[11'h017] = 8'h69;
    mem[11'h018] = 8'ha2;
    mem[11'h019] = 8'h6f;
    mem[11'h01a] = 8'h9d;
    mem[11'h01b] = 8'h73;
    mem[11'h01c] = 8'h99;
    mem[11'h01d] = 8'h77;
    mem[11'h01e] = 8'h95;
    mem[11'h01f] = 8'h7b;
    mem[11'h020] = 8'h91;
    mem[11'h021] = 8'h7f;
    mem[11'h022] = 8'h8e;
    mem[11'h023] = 8'h82;
    mem[11'h024] = 8'h8a;
    mem[11'h025] = 8'h85;
    mem[11'h026] = 8'h87;
    mem[11'h027] = 8'h89;
    mem[11'h028] = 8'h84;
    mem[11'h029] = 8'h8c;
    mem[11'h02a] = 8'h80;
    mem[11'h02b] = 8'h8f;
    mem[11'h02c] = 8'h7d;
    mem[11'h02d] = 8'h3c;
    mem[11'h02e] = 8'h19;
    mem[11'h02f] = 8'h3c;
    mem[11'h030] = 8'h7a;
    mem[11'h031] = 8'h37;
    mem[11'h032] = 8'h25;
    mem[11'h033] = 8'h37;
    mem[11'h034] = 8'h77;
    mem[11'h035] = 8'h34;
    mem[11'h036] = 8'h2f;
    mem[11'h037] = 8'h34;
    mem[11'h038] = 8'h74;
    mem[11'h039] = 8'h31;
    mem[11'h03a] = 8'h38;
    mem[11'h03b] = 8'h30;
    mem[11'h03c] = 8'h72;
    mem[11'h03d] = 8'h2e;
    mem[11'h03e] = 8'h3f;
    mem[11'h03f] = 8'h2e;
    mem[11'h040] = 8'h6f;
    mem[11'h041] = 8'h2d;
    mem[11'h042] = 8'h45;
    mem[11'h043] = 8'h2d;
    mem[11'h044] = 8'h6c;
    mem[11'h045] = 8'h2b;
    mem[11'h046] = 8'h4b;
    mem[11'h047] = 8'h2b;
    mem[11'h048] = 8'h6a;
    mem[11'h049] = 8'h29;
    mem[11'h04a] = 8'h51;
    mem[11'h04b] = 8'h29;
    mem[11'h04c] = 8'h68;
    mem[11'h04d] = 8'h28;
    mem[11'h04e] = 8'h55;
    mem[11'h04f] = 8'h29;
    mem[11'h050] = 8'h64;
    mem[11'h051] = 8'h28;
    mem[11'h052] = 8'h59;
    mem[11'h053] = 8'h28;
    mem[11'h054] = 8'h62;
    mem[11'h055] = 8'h27;
    mem[11'h056] = 8'h5e;
    mem[11'h057] = 8'h26;
    mem[11'h058] = 8'h60;
    mem[11'h059] = 8'h25;
    mem[11'h05a] = 8'h63;
    mem[11'h05b] = 8'h25;
    mem[11'h05c] = 8'h5e;
    mem[11'h05d] = 8'h24;
    mem[11'h05e] = 8'h67;
    mem[11'h05f] = 8'h24;
    mem[11'h060] = 8'h5c;
    mem[11'h061] = 8'h24;
    mem[11'h062] = 8'h6a;
    mem[11'h063] = 8'h23;
    mem[11'h064] = 8'h5a;
    mem[11'h065] = 8'h23;
    mem[11'h066] = 8'h6d;
    mem[11'h067] = 8'h23;
    mem[11'h068] = 8'h58;
    mem[11'h069] = 8'h22;
    mem[11'h06a] = 8'h71;
    mem[11'h06b] = 8'h23;
    mem[11'h06c] = 8'h55;
    mem[11'h06d] = 8'h21;
    mem[11'h06e] = 8'h75;
    mem[11'h06f] = 8'h22;
    mem[11'h070] = 8'h53;
    mem[11'h071] = 8'h21;
    mem[11'h072] = 8'h77;
    mem[11'h073] = 8'h22;
    mem[11'h074] = 8'h51;
    mem[11'h075] = 8'h20;
    mem[11'h076] = 8'h7b;
    mem[11'h077] = 8'h21;
    mem[11'h078] = 8'h4f;
    mem[11'h079] = 8'h20;
    mem[11'h07a] = 8'h7d;
    mem[11'h07b] = 8'h21;
    mem[11'h07c] = 8'h4d;
    mem[11'h07d] = 8'h1f;
    mem[11'h07e] = 8'h81;
    mem[11'h07f] = 8'h1f;
    mem[11'h080] = 8'h4c;
    mem[11'h081] = 8'h1f;
    mem[11'h082] = 8'h83;
    mem[11'h083] = 8'h1f;
    mem[11'h084] = 8'h4a;
    mem[11'h085] = 8'h1f;
    mem[11'h086] = 8'h85;
    mem[11'h087] = 8'h1f;
    mem[11'h088] = 8'h48;
    mem[11'h089] = 8'h1e;
    mem[11'h08a] = 8'h89;
    mem[11'h08b] = 8'h1e;
    mem[11'h08c] = 8'h46;
    mem[11'h08d] = 8'h1e;
    mem[11'h08e] = 8'h8b;
    mem[11'h08f] = 8'h1e;
    mem[11'h090] = 8'h44;
    mem[11'h091] = 8'h1e;
    mem[11'h092] = 8'h8d;
    mem[11'h093] = 8'h1e;
    mem[11'h094] = 8'h42;
    mem[11'h095] = 8'h1e;
    mem[11'h096] = 8'h8f;
    mem[11'h097] = 8'h1e;
    mem[11'h098] = 8'h40;
    mem[11'h099] = 8'h1d;
    mem[11'h09a] = 8'h93;
    mem[11'h09b] = 8'h1d;
    mem[11'h09c] = 8'h3f;
    mem[11'h09d] = 8'h1c;
    mem[11'h09e] = 8'h95;
    mem[11'h09f] = 8'h1c;
    mem[11'h0a0] = 8'h3e;
    mem[11'h0a1] = 8'h1c;
    mem[11'h0a2] = 8'h97;
    mem[11'h0a3] = 8'h1c;
    mem[11'h0a4] = 8'h3c;
    mem[11'h0a5] = 8'h1c;
    mem[11'h0a6] = 8'h99;
    mem[11'h0a7] = 8'h1c;
    mem[11'h0a8] = 8'h3a;
    mem[11'h0a9] = 8'h1c;
    mem[11'h0aa] = 8'h9b;
    mem[11'h0ab] = 8'h1c;
    mem[11'h0ac] = 8'h39;
    mem[11'h0ad] = 8'h1b;
    mem[11'h0ae] = 8'h9d;
    mem[11'h0af] = 8'h1c;
    mem[11'h0b0] = 8'h37;
    mem[11'h0b1] = 8'h1b;
    mem[11'h0b2] = 8'h9f;
    mem[11'h0b3] = 8'h1b;
    mem[11'h0b4] = 8'h36;
    mem[11'h0b5] = 8'h86;
    mem[11'h0b6] = 8'h36;
    mem[11'h0b7] = 8'h1b;
    mem[11'h0b8] = 8'h34;
    mem[11'h0b9] = 8'h87;
    mem[11'h0ba] = 8'h37;
    mem[11'h0bb] = 8'h1b;
    mem[11'h0bc] = 8'h33;
    mem[11'h0bd] = 8'h87;
    mem[11'h0be] = 8'h38;
    mem[11'h0bf] = 8'h1a;
    mem[11'h0c0] = 8'h32;
    mem[11'h0c1] = 8'h88;
    mem[11'h0c2] = 8'h39;
    mem[11'h0c3] = 8'h1a;
    mem[11'h0c4] = 8'h30;
    mem[11'h0c5] = 8'h89;
    mem[11'h0c6] = 8'h3a;
    mem[11'h0c7] = 8'h1a;
    mem[11'h0c8] = 8'h2f;
    mem[11'h0c9] = 8'h89;
    mem[11'h0ca] = 8'h3a;
    mem[11'h0cb] = 8'h1a;
    mem[11'h0cc] = 8'h2e;
    mem[11'h0cd] = 8'h8a;
    mem[11'h0ce] = 8'h3b;
    mem[11'h0cf] = 8'h1a;
    mem[11'h0d0] = 8'h2c;
    mem[11'h0d1] = 8'h8b;
    mem[11'h0d2] = 8'h3c;
    mem[11'h0d3] = 8'h1a;
    mem[11'h0d4] = 8'h2b;
    mem[11'h0d5] = 8'h8b;
    mem[11'h0d6] = 8'h3d;
    mem[11'h0d7] = 8'h19;
    mem[11'h0d8] = 8'h2a;
    mem[11'h0d9] = 8'h8c;
    mem[11'h0da] = 8'h3e;
    mem[11'h0db] = 8'h19;
    mem[11'h0dc] = 8'h29;
    mem[11'h0dd] = 8'h8c;
    mem[11'h0de] = 8'h3e;
    mem[11'h0df] = 8'h19;
    mem[11'h0e0] = 8'h28;
    mem[11'h0e1] = 8'h8d;
    mem[11'h0e2] = 8'h3f;
    mem[11'h0e3] = 8'h19;
    mem[11'h0e4] = 8'h27;
    mem[11'h0e5] = 8'h8d;
    mem[11'h0e6] = 8'h40;
    mem[11'h0e7] = 8'h19;
    mem[11'h0e8] = 8'h25;
    mem[11'h0e9] = 8'h8e;
    mem[11'h0ea] = 8'h41;
    mem[11'h0eb] = 8'h18;
    mem[11'h0ec] = 8'h24;
    mem[11'h0ed] = 8'h8f;
    mem[11'h0ee] = 8'h41;
    mem[11'h0ef] = 8'h19;
    mem[11'h0f0] = 8'h23;
    mem[11'h0f1] = 8'h8f;
    mem[11'h0f2] = 8'h42;
    mem[11'h0f3] = 8'h18;
    mem[11'h0f4] = 8'h22;
    mem[11'h0f5] = 8'h90;
    mem[11'h0f6] = 8'h43;
    mem[11'h0f7] = 8'h18;
    mem[11'h0f8] = 8'h21;
    mem[11'h0f9] = 8'h90;
    mem[11'h0fa] = 8'h43;
    mem[11'h0fb] = 8'h18;
    mem[11'h0fc] = 8'h20;
    mem[11'h0fd] = 8'h91;
    mem[11'h0fe] = 8'h44;
    mem[11'h0ff] = 8'h18;
    mem[11'h100] = 8'h1f;
    mem[11'h101] = 8'h91;
    mem[11'h102] = 8'h45;
    mem[11'h103] = 8'h17;
    mem[11'h104] = 8'h1e;
    mem[11'h105] = 8'h92;
    mem[11'h106] = 8'h45;
    mem[11'h107] = 8'h18;
    mem[11'h108] = 8'h1d;
    mem[11'h109] = 8'h92;
    mem[11'h10a] = 8'h46;
    mem[11'h10b] = 8'h17;
    mem[11'h10c] = 8'h1c;
    mem[11'h10d] = 8'h93;
    mem[11'h10e] = 8'h46;
    mem[11'h10f] = 8'h18;
    mem[11'h110] = 8'h1b;
    mem[11'h111] = 8'h93;
    mem[11'h112] = 8'h47;
    mem[11'h113] = 8'h17;
    mem[11'h114] = 8'h1b;
    mem[11'h115] = 8'h93;
    mem[11'h116] = 8'h48;
    mem[11'h117] = 8'h17;
    mem[11'h118] = 8'h19;
    mem[11'h119] = 8'h94;
    mem[11'h11a] = 8'h48;
    mem[11'h11b] = 8'h17;
    mem[11'h11c] = 8'h19;
    mem[11'h11d] = 8'h94;
    mem[11'h11e] = 8'h49;
    mem[11'h11f] = 8'h16;
    mem[11'h120] = 8'h18;
    mem[11'h121] = 8'h95;
    mem[11'h122] = 8'h49;
    mem[11'h123] = 8'h17;
    mem[11'h124] = 8'h17;
    mem[11'h125] = 8'h95;
    mem[11'h126] = 8'h4a;
    mem[11'h127] = 8'h16;
    mem[11'h128] = 8'h16;
    mem[11'h129] = 8'h96;
    mem[11'h12a] = 8'h4a;
    mem[11'h12b] = 8'h17;
    mem[11'h12c] = 8'h15;
    mem[11'h12d] = 8'h96;
    mem[11'h12e] = 8'h4b;
    mem[11'h12f] = 8'h16;
    mem[11'h130] = 8'h15;
    mem[11'h131] = 8'h96;
    mem[11'h132] = 8'h4b;
    mem[11'h133] = 8'h16;
    mem[11'h134] = 8'h14;
    mem[11'h135] = 8'h97;
    mem[11'h136] = 8'h4c;
    mem[11'h137] = 8'h16;
    mem[11'h138] = 8'h13;
    mem[11'h139] = 8'h97;
    mem[11'h13a] = 8'h4c;
    mem[11'h13b] = 8'h16;
    mem[11'h13c] = 8'h13;
    mem[11'h13d] = 8'h97;
    mem[11'h13e] = 8'h4c;
    mem[11'h13f] = 8'h16;
    mem[11'h140] = 8'h12;
    mem[11'h141] = 8'h98;
    mem[11'h142] = 8'h4d;
    mem[11'h143] = 8'h16;
    mem[11'h144] = 8'h11;
    mem[11'h145] = 8'h98;
    mem[11'h146] = 8'h4d;
    mem[11'h147] = 8'h16;
    mem[11'h148] = 8'h5b;
    mem[11'h149] = 8'h27;
    mem[11'h14a] = 8'h75;
    mem[11'h14b] = 8'h16;
    mem[11'h14c] = 8'h5a;
    mem[11'h14d] = 8'h27;
    mem[11'h14e] = 8'h75;
    mem[11'h14f] = 8'h16;
    mem[11'h150] = 8'h5a;
    mem[11'h151] = 8'h27;
    mem[11'h152] = 8'h75;
    mem[11'h153] = 8'h16;
    mem[11'h154] = 8'h5a;
    mem[11'h155] = 8'h27;
    mem[11'h156] = 8'h76;
    mem[11'h157] = 8'h15;
    mem[11'h158] = 8'h5a;
    mem[11'h159] = 8'h27;
    mem[11'h15a] = 8'h76;
    mem[11'h15b] = 8'h16;
    mem[11'h15c] = 8'h59;
    mem[11'h15d] = 8'h27;
    mem[11'h15e] = 8'h76;
    mem[11'h15f] = 8'h16;
    mem[11'h160] = 8'h59;
    mem[11'h161] = 8'h27;
    mem[11'h162] = 8'h77;
    mem[11'h163] = 8'h15;
    mem[11'h164] = 8'h59;
    mem[11'h165] = 8'h27;
    mem[11'h166] = 8'h77;
    mem[11'h167] = 8'h16;
    mem[11'h168] = 8'h58;
    mem[11'h169] = 8'h27;
    mem[11'h16a] = 8'h77;
    mem[11'h16b] = 8'h16;
    mem[11'h16c] = 8'h58;
    mem[11'h16d] = 8'h27;
    mem[11'h16e] = 8'h78;
    mem[11'h16f] = 8'h15;
    mem[11'h170] = 8'h58;
    mem[11'h171] = 8'h27;
    mem[11'h172] = 8'h78;
    mem[11'h173] = 8'h15;
    mem[11'h174] = 8'h0b;
    mem[11'h175] = 8'h15;
    mem[11'h176] = 8'h36;
    mem[11'h177] = 8'h27;
    mem[11'h178] = 8'h78;
    mem[11'h179] = 8'h15;
    mem[11'h17a] = 8'h0a;
    mem[11'h17b] = 8'h16;
    mem[11'h17c] = 8'h36;
    mem[11'h17d] = 8'h27;
    mem[11'h17e] = 8'h79;
    mem[11'h17f] = 8'h15;
    mem[11'h180] = 8'h09;
    mem[11'h181] = 8'h15;
    mem[11'h182] = 8'h37;
    mem[11'h183] = 8'h27;
    mem[11'h184] = 8'h79;
    mem[11'h185] = 8'h15;
    mem[11'h186] = 8'h09;
    mem[11'h187] = 8'h15;
    mem[11'h188] = 8'h37;
    mem[11'h189] = 8'h27;
    mem[11'h18a] = 8'h79;
    mem[11'h18b] = 8'h15;
    mem[11'h18c] = 8'h09;
    mem[11'h18d] = 8'h15;
    mem[11'h18e] = 8'h37;
    mem[11'h18f] = 8'h27;
    mem[11'h190] = 8'h79;
    mem[11'h191] = 8'h15;
    mem[11'h192] = 8'h09;
    mem[11'h193] = 8'h15;
    mem[11'h194] = 8'h37;
    mem[11'h195] = 8'h27;
    mem[11'h196] = 8'h7a;
    mem[11'h197] = 8'h14;
    mem[11'h198] = 8'h08;
    mem[11'h199] = 8'h15;
    mem[11'h19a] = 8'h38;
    mem[11'h19b] = 8'h27;
    mem[11'h19c] = 8'h7a;
    mem[11'h19d] = 8'h15;
    mem[11'h19e] = 8'h07;
    mem[11'h19f] = 8'h15;
    mem[11'h1a0] = 8'h38;
    mem[11'h1a1] = 8'h27;
    mem[11'h1a2] = 8'h7a;
    mem[11'h1a3] = 8'h15;
    mem[11'h1a4] = 8'h07;
    mem[11'h1a5] = 8'h15;
    mem[11'h1a6] = 8'h38;
    mem[11'h1a7] = 8'h27;
    mem[11'h1a8] = 8'h7a;
    mem[11'h1a9] = 8'h15;
    mem[11'h1aa] = 8'h07;
    mem[11'h1ab] = 8'h15;
    mem[11'h1ac] = 8'h38;
    mem[11'h1ad] = 8'h27;
    mem[11'h1ae] = 8'h7a;
    mem[11'h1af] = 8'h15;
    mem[11'h1b0] = 8'h07;
    mem[11'h1b1] = 8'h15;
    mem[11'h1b2] = 8'h38;
    mem[11'h1b3] = 8'h27;
    mem[11'h1b4] = 8'h7b;
    mem[11'h1b5] = 8'h14;
    mem[11'h1b6] = 8'h07;
    mem[11'h1b7] = 8'h14;
    mem[11'h1b8] = 8'h39;
    mem[11'h1b9] = 8'h27;
    mem[11'h1ba] = 8'h7b;
    mem[11'h1bb] = 8'h14;
    mem[11'h1bc] = 8'h06;
    mem[11'h1bd] = 8'h15;
    mem[11'h1be] = 8'h39;
    mem[11'h1bf] = 8'h27;
    mem[11'h1c0] = 8'h7b;
    mem[11'h1c1] = 8'h15;
    mem[11'h1c2] = 8'h05;
    mem[11'h1c3] = 8'h15;
    mem[11'h1c4] = 8'h39;
    mem[11'h1c5] = 8'h27;
    mem[11'h1c6] = 8'h7b;
    mem[11'h1c7] = 8'h15;
    mem[11'h1c8] = 8'h05;
    mem[11'h1c9] = 8'h15;
    mem[11'h1ca] = 8'h39;
    mem[11'h1cb] = 8'h27;
    mem[11'h1cc] = 8'h7b;
    mem[11'h1cd] = 8'h15;
    mem[11'h1ce] = 8'h05;
    mem[11'h1cf] = 8'h15;
    mem[11'h1d0] = 8'h39;
    mem[11'h1d1] = 8'h27;
    mem[11'h1d2] = 8'h7b;
    mem[11'h1d3] = 8'h15;
    mem[11'h1d4] = 8'h05;
    mem[11'h1d5] = 8'h15;
    mem[11'h1d6] = 8'h39;
    mem[11'h1d7] = 8'h27;
    mem[11'h1d8] = 8'h7b;
    mem[11'h1d9] = 8'h15;
    mem[11'h1da] = 8'h05;
    mem[11'h1db] = 8'h14;
    mem[11'h1dc] = 8'h3a;
    mem[11'h1dd] = 8'h27;
    mem[11'h1de] = 8'h7c;
    mem[11'h1df] = 8'h14;
    mem[11'h1e0] = 8'h05;
    mem[11'h1e1] = 8'h14;
    mem[11'h1e2] = 8'h3a;
    mem[11'h1e3] = 8'h8c;
    mem[11'h1e4] = 8'h17;
    mem[11'h1e5] = 8'h14;
    mem[11'h1e6] = 8'h05;
    mem[11'h1e7] = 8'h14;
    mem[11'h1e8] = 8'h3a;
    mem[11'h1e9] = 8'h8c;
    mem[11'h1ea] = 8'h17;
    mem[11'h1eb] = 8'h14;
    mem[11'h1ec] = 8'h05;
    mem[11'h1ed] = 8'h14;
    mem[11'h1ee] = 8'h3a;
    mem[11'h1ef] = 8'h8c;
    mem[11'h1f0] = 8'h17;
    mem[11'h1f1] = 8'h14;
    mem[11'h1f2] = 8'h05;
    mem[11'h1f3] = 8'h14;
    mem[11'h1f4] = 8'h3a;
    mem[11'h1f5] = 8'h8c;
    mem[11'h1f6] = 8'h17;
    mem[11'h1f7] = 8'h14;
    mem[11'h1f8] = 8'h05;
    mem[11'h1f9] = 8'h14;
    mem[11'h1fa] = 8'h3a;
    mem[11'h1fb] = 8'h8c;
    mem[11'h1fc] = 8'h17;
    mem[11'h1fd] = 8'h15;
    mem[11'h1fe] = 8'h04;
    mem[11'h1ff] = 8'h14;
    mem[11'h200] = 8'h3a;
    mem[11'h201] = 8'h8c;
    mem[11'h202] = 8'h17;
    mem[11'h203] = 8'h15;
    mem[11'h204] = 8'h04;
    mem[11'h205] = 8'h14;
    mem[11'h206] = 8'h3a;
    mem[11'h207] = 8'h8c;
    mem[11'h208] = 8'h17;
    mem[11'h209] = 8'h15;
    mem[11'h20a] = 8'h03;
    mem[11'h20b] = 8'h15;
    mem[11'h20c] = 8'h3a;
    mem[11'h20d] = 8'h8c;
    mem[11'h20e] = 8'h17;
    mem[11'h20f] = 8'h15;
    mem[11'h210] = 8'h03;
    mem[11'h211] = 8'h15;
    mem[11'h212] = 8'h3a;
    mem[11'h213] = 8'h8c;
    mem[11'h214] = 8'h17;
    mem[11'h215] = 8'h15;
    mem[11'h216] = 8'h03;
    mem[11'h217] = 8'h15;
    mem[11'h218] = 8'h3a;
    mem[11'h219] = 8'h8c;
    mem[11'h21a] = 8'h17;
    mem[11'h21b] = 8'h15;
    mem[11'h21c] = 8'h03;
    mem[11'h21d] = 8'h15;
    mem[11'h21e] = 8'h3a;
    mem[11'h21f] = 8'h8c;
    mem[11'h220] = 8'h17;
    mem[11'h221] = 8'h15;
    mem[11'h222] = 8'h03;
    mem[11'h223] = 8'h15;
    mem[11'h224] = 8'h3a;
    mem[11'h225] = 8'h8c;
    mem[11'h226] = 8'h17;
    mem[11'h227] = 8'h15;
    mem[11'h228] = 8'h03;
    mem[11'h229] = 8'h15;
    mem[11'h22a] = 8'h3a;
    mem[11'h22b] = 8'h8c;
    mem[11'h22c] = 8'h17;
    mem[11'h22d] = 8'h15;
    mem[11'h22e] = 8'h03;
    mem[11'h22f] = 8'h15;
    mem[11'h230] = 8'h3a;
    mem[11'h231] = 8'h8c;
    mem[11'h232] = 8'h17;
    mem[11'h233] = 8'h15;
    mem[11'h234] = 8'h03;
    mem[11'h235] = 8'h15;
    mem[11'h236] = 8'h3a;
    mem[11'h237] = 8'h8c;
    mem[11'h238] = 8'h17;
    mem[11'h239] = 8'h15;
    mem[11'h23a] = 8'h03;
    mem[11'h23b] = 8'h15;
    mem[11'h23c] = 8'h3a;
    mem[11'h23d] = 8'h8c;
    mem[11'h23e] = 8'h17;
    mem[11'h23f] = 8'h15;
    mem[11'h240] = 8'h03;
    mem[11'h241] = 8'h15;
    mem[11'h242] = 8'h3a;
    mem[11'h243] = 8'h8c;
    mem[11'h244] = 8'h17;
    mem[11'h245] = 8'h15;
    mem[11'h246] = 8'h03;
    mem[11'h247] = 8'h15;
    mem[11'h248] = 8'h3a;
    mem[11'h249] = 8'h8c;
    mem[11'h24a] = 8'h17;
    mem[11'h24b] = 8'h15;
    mem[11'h24c] = 8'h04;
    mem[11'h24d] = 8'h14;
    mem[11'h24e] = 8'h3a;
    mem[11'h24f] = 8'h8c;
    mem[11'h250] = 8'h17;
    mem[11'h251] = 8'h15;
    mem[11'h252] = 8'h04;
    mem[11'h253] = 8'h14;
    mem[11'h254] = 8'h3a;
    mem[11'h255] = 8'h8c;
    mem[11'h256] = 8'h17;
    mem[11'h257] = 8'h15;
    mem[11'h258] = 8'h04;
    mem[11'h259] = 8'h14;
    mem[11'h25a] = 8'h3a;
    mem[11'h25b] = 8'h8c;
    mem[11'h25c] = 8'h17;
    mem[11'h25d] = 8'h14;
    mem[11'h25e] = 8'h05;
    mem[11'h25f] = 8'h14;
    mem[11'h260] = 8'h3a;
    mem[11'h261] = 8'h8c;
    mem[11'h262] = 8'h17;
    mem[11'h263] = 8'h14;
    mem[11'h264] = 8'h05;
    mem[11'h265] = 8'h14;
    mem[11'h266] = 8'h3a;
    mem[11'h267] = 8'h8c;
    mem[11'h268] = 8'h17;
    mem[11'h269] = 8'h14;
    mem[11'h26a] = 8'h05;
    mem[11'h26b] = 8'h14;
    mem[11'h26c] = 8'h3a;
    mem[11'h26d] = 8'h8c;
    mem[11'h26e] = 8'h17;
    mem[11'h26f] = 8'h14;
    mem[11'h270] = 8'h05;
    mem[11'h271] = 8'h14;
    mem[11'h272] = 8'h3a;
    mem[11'h273] = 8'h8c;
    mem[11'h274] = 8'h17;
    mem[11'h275] = 8'h14;
    mem[11'h276] = 8'h05;
    mem[11'h277] = 8'h15;
    mem[11'h278] = 8'h39;
    mem[11'h279] = 8'h8c;
    mem[11'h27a] = 8'h17;
    mem[11'h27b] = 8'h14;
    mem[11'h27c] = 8'h05;
    mem[11'h27d] = 8'h15;
    mem[11'h27e] = 8'h39;
    mem[11'h27f] = 8'h8c;
    mem[11'h280] = 8'h16;
    mem[11'h281] = 8'h15;
    mem[11'h282] = 8'h05;
    mem[11'h283] = 8'h15;
    mem[11'h284] = 8'h39;
    mem[11'h285] = 8'h8c;
    mem[11'h286] = 8'h16;
    mem[11'h287] = 8'h15;
    mem[11'h288] = 8'h05;
    mem[11'h289] = 8'h15;
    mem[11'h28a] = 8'h39;
    mem[11'h28b] = 8'h8c;
    mem[11'h28c] = 8'h16;
    mem[11'h28d] = 8'h15;
    mem[11'h28e] = 8'h05;
    mem[11'h28f] = 8'h15;
    mem[11'h290] = 8'h39;
    mem[11'h291] = 8'h8c;
    mem[11'h292] = 8'h16;
    mem[11'h293] = 8'h15;
    mem[11'h294] = 8'h06;
    mem[11'h295] = 8'h14;
    mem[11'h296] = 8'h39;
    mem[11'h297] = 8'h8c;
    mem[11'h298] = 8'h16;
    mem[11'h299] = 8'h15;
    mem[11'h29a] = 8'h06;
    mem[11'h29b] = 8'h14;
    mem[11'h29c] = 8'h39;
    mem[11'h29d] = 8'h8c;
    mem[11'h29e] = 8'h16;
    mem[11'h29f] = 8'h14;
    mem[11'h2a0] = 8'h07;
    mem[11'h2a1] = 8'h15;
    mem[11'h2a2] = 8'h38;
    mem[11'h2a3] = 8'h8c;
    mem[11'h2a4] = 8'h15;
    mem[11'h2a5] = 8'h15;
    mem[11'h2a6] = 8'h07;
    mem[11'h2a7] = 8'h15;
    mem[11'h2a8] = 8'h38;
    mem[11'h2a9] = 8'h8c;
    mem[11'h2aa] = 8'h15;
    mem[11'h2ab] = 8'h15;
    mem[11'h2ac] = 8'h07;
    mem[11'h2ad] = 8'h15;
    mem[11'h2ae] = 8'h38;
    mem[11'h2af] = 8'h8c;
    mem[11'h2b0] = 8'h15;
    mem[11'h2b1] = 8'h15;
    mem[11'h2b2] = 8'h07;
    mem[11'h2b3] = 8'h15;
    mem[11'h2b4] = 8'h38;
    mem[11'h2b5] = 8'h8c;
    mem[11'h2b6] = 8'h15;
    mem[11'h2b7] = 8'h15;
    mem[11'h2b8] = 8'h08;
    mem[11'h2b9] = 8'h14;
    mem[11'h2ba] = 8'h38;
    mem[11'h2bb] = 8'h8c;
    mem[11'h2bc] = 8'h15;
    mem[11'h2bd] = 8'h15;
    mem[11'h2be] = 8'h08;
    mem[11'h2bf] = 8'h15;
    mem[11'h2c0] = 8'h37;
    mem[11'h2c1] = 8'h27;
    mem[11'h2c2] = 8'h15;
    mem[11'h2c3] = 8'h27;
    mem[11'h2c4] = 8'h3b;
    mem[11'h2c5] = 8'h15;
    mem[11'h2c6] = 8'h09;
    mem[11'h2c7] = 8'h15;
    mem[11'h2c8] = 8'h37;
    mem[11'h2c9] = 8'h27;
    mem[11'h2ca] = 8'h15;
    mem[11'h2cb] = 8'h27;
    mem[11'h2cc] = 8'h3b;
    mem[11'h2cd] = 8'h15;
    mem[11'h2ce] = 8'h09;
    mem[11'h2cf] = 8'h15;
    mem[11'h2d0] = 8'h37;
    mem[11'h2d1] = 8'h27;
    mem[11'h2d2] = 8'h15;
    mem[11'h2d3] = 8'h27;
    mem[11'h2d4] = 8'h3b;
    mem[11'h2d5] = 8'h15;
    mem[11'h2d6] = 8'h09;
    mem[11'h2d7] = 8'h15;
    mem[11'h2d8] = 8'h37;
    mem[11'h2d9] = 8'h27;
    mem[11'h2da] = 8'h15;
    mem[11'h2db] = 8'h27;
    mem[11'h2dc] = 8'h3b;
    mem[11'h2dd] = 8'h15;
    mem[11'h2de] = 8'h0a;
    mem[11'h2df] = 8'h15;
    mem[11'h2e0] = 8'h36;
    mem[11'h2e1] = 8'h27;
    mem[11'h2e2] = 8'h15;
    mem[11'h2e3] = 8'h27;
    mem[11'h2e4] = 8'h3a;
    mem[11'h2e5] = 8'h16;
    mem[11'h2e6] = 8'h0a;
    mem[11'h2e7] = 8'h15;
    mem[11'h2e8] = 8'h36;
    mem[11'h2e9] = 8'h27;
    mem[11'h2ea] = 8'h15;
    mem[11'h2eb] = 8'h27;
    mem[11'h2ec] = 8'h3a;
    mem[11'h2ed] = 8'h15;
    mem[11'h2ee] = 8'h0b;
    mem[11'h2ef] = 8'h15;
    mem[11'h2f0] = 8'h36;
    mem[11'h2f1] = 8'h27;
    mem[11'h2f2] = 8'h15;
    mem[11'h2f3] = 8'h27;
    mem[11'h2f4] = 8'h3a;
    mem[11'h2f5] = 8'h15;
    mem[11'h2f6] = 8'h0b;
    mem[11'h2f7] = 8'h16;
    mem[11'h2f8] = 8'h35;
    mem[11'h2f9] = 8'h27;
    mem[11'h2fa] = 8'h15;
    mem[11'h2fb] = 8'h27;
    mem[11'h2fc] = 8'h39;
    mem[11'h2fd] = 8'h16;
    mem[11'h2fe] = 8'h0c;
    mem[11'h2ff] = 8'h15;
    mem[11'h300] = 8'h35;
    mem[11'h301] = 8'h27;
    mem[11'h302] = 8'h15;
    mem[11'h303] = 8'h27;
    mem[11'h304] = 8'h39;
    mem[11'h305] = 8'h16;
    mem[11'h306] = 8'h0c;
    mem[11'h307] = 8'h15;
    mem[11'h308] = 8'h35;
    mem[11'h309] = 8'h27;
    mem[11'h30a] = 8'h15;
    mem[11'h30b] = 8'h27;
    mem[11'h30c] = 8'h39;
    mem[11'h30d] = 8'h15;
    mem[11'h30e] = 8'h0d;
    mem[11'h30f] = 8'h16;
    mem[11'h310] = 8'h34;
    mem[11'h311] = 8'h27;
    mem[11'h312] = 8'h15;
    mem[11'h313] = 8'h27;
    mem[11'h314] = 8'h39;
    mem[11'h315] = 8'h15;
    mem[11'h316] = 8'h0d;
    mem[11'h317] = 8'h16;
    mem[11'h318] = 8'h34;
    mem[11'h319] = 8'h27;
    mem[11'h31a] = 8'h15;
    mem[11'h31b] = 8'h27;
    mem[11'h31c] = 8'h38;
    mem[11'h31d] = 8'h16;
    mem[11'h31e] = 8'h0e;
    mem[11'h31f] = 8'h15;
    mem[11'h320] = 8'h34;
    mem[11'h321] = 8'h27;
    mem[11'h322] = 8'h15;
    mem[11'h323] = 8'h27;
    mem[11'h324] = 8'h38;
    mem[11'h325] = 8'h16;
    mem[11'h326] = 8'h0e;
    mem[11'h327] = 8'h16;
    mem[11'h328] = 8'h33;
    mem[11'h329] = 8'h27;
    mem[11'h32a] = 8'h15;
    mem[11'h32b] = 8'h27;
    mem[11'h32c] = 8'h37;
    mem[11'h32d] = 8'h16;
    mem[11'h32e] = 8'h0f;
    mem[11'h32f] = 8'h16;
    mem[11'h330] = 8'h33;
    mem[11'h331] = 8'h27;
    mem[11'h332] = 8'h15;
    mem[11'h333] = 8'h27;
    mem[11'h334] = 8'h37;
    mem[11'h335] = 8'h16;
    mem[11'h336] = 8'h10;
    mem[11'h337] = 8'h15;
    mem[11'h338] = 8'h33;
    mem[11'h339] = 8'h27;
    mem[11'h33a] = 8'h15;
    mem[11'h33b] = 8'h27;
    mem[11'h33c] = 8'h37;
    mem[11'h33d] = 8'h16;
    mem[11'h33e] = 8'h10;
    mem[11'h33f] = 8'h16;
    mem[11'h340] = 8'h32;
    mem[11'h341] = 8'h27;
    mem[11'h342] = 8'h15;
    mem[11'h343] = 8'h27;
    mem[11'h344] = 8'h36;
    mem[11'h345] = 8'h16;
    mem[11'h346] = 8'h11;
    mem[11'h347] = 8'h16;
    mem[11'h348] = 8'h32;
    mem[11'h349] = 8'h27;
    mem[11'h34a] = 8'h15;
    mem[11'h34b] = 8'h27;
    mem[11'h34c] = 8'h36;
    mem[11'h34d] = 8'h16;
    mem[11'h34e] = 8'h12;
    mem[11'h34f] = 8'h16;
    mem[11'h350] = 8'h31;
    mem[11'h351] = 8'h27;
    mem[11'h352] = 8'h15;
    mem[11'h353] = 8'h27;
    mem[11'h354] = 8'h35;
    mem[11'h355] = 8'h17;
    mem[11'h356] = 8'h12;
    mem[11'h357] = 8'h16;
    mem[11'h358] = 8'h31;
    mem[11'h359] = 8'h27;
    mem[11'h35a] = 8'h15;
    mem[11'h35b] = 8'h27;
    mem[11'h35c] = 8'h35;
    mem[11'h35d] = 8'h16;
    mem[11'h35e] = 8'h13;
    mem[11'h35f] = 8'h16;
    mem[11'h360] = 8'h31;
    mem[11'h361] = 8'h27;
    mem[11'h362] = 8'h15;
    mem[11'h363] = 8'h27;
    mem[11'h364] = 8'h35;
    mem[11'h365] = 8'h16;
    mem[11'h366] = 8'h14;
    mem[11'h367] = 8'h16;
    mem[11'h368] = 8'h30;
    mem[11'h369] = 8'h27;
    mem[11'h36a] = 8'h15;
    mem[11'h36b] = 8'h27;
    mem[11'h36c] = 8'h34;
    mem[11'h36d] = 8'h17;
    mem[11'h36e] = 8'h14;
    mem[11'h36f] = 8'h16;
    mem[11'h370] = 8'h30;
    mem[11'h371] = 8'h27;
    mem[11'h372] = 8'h15;
    mem[11'h373] = 8'h27;
    mem[11'h374] = 8'h34;
    mem[11'h375] = 8'h16;
    mem[11'h376] = 8'h15;
    mem[11'h377] = 8'h17;
    mem[11'h378] = 8'h2f;
    mem[11'h379] = 8'h27;
    mem[11'h37a] = 8'h15;
    mem[11'h37b] = 8'h27;
    mem[11'h37c] = 8'h33;
    mem[11'h37d] = 8'h17;
    mem[11'h37e] = 8'h16;
    mem[11'h37f] = 8'h16;
    mem[11'h380] = 8'h6d;
    mem[11'h381] = 8'h27;
    mem[11'h382] = 8'h33;
    mem[11'h383] = 8'h16;
    mem[11'h384] = 8'h17;
    mem[11'h385] = 8'h17;
    mem[11'h386] = 8'h6c;
    mem[11'h387] = 8'h27;
    mem[11'h388] = 8'h32;
    mem[11'h389] = 8'h17;
    mem[11'h38a] = 8'h18;
    mem[11'h38b] = 8'h16;
    mem[11'h38c] = 8'h6c;
    mem[11'h38d] = 8'h27;
    mem[11'h38e] = 8'h32;
    mem[11'h38f] = 8'h17;
    mem[11'h390] = 8'h18;
    mem[11'h391] = 8'h17;
    mem[11'h392] = 8'h6b;
    mem[11'h393] = 8'h27;
    mem[11'h394] = 8'h31;
    mem[11'h395] = 8'h17;
    mem[11'h396] = 8'h19;
    mem[11'h397] = 8'h17;
    mem[11'h398] = 8'h6b;
    mem[11'h399] = 8'h27;
    mem[11'h39a] = 8'h31;
    mem[11'h39b] = 8'h17;
    mem[11'h39c] = 8'h1a;
    mem[11'h39d] = 8'h17;
    mem[11'h39e] = 8'h6a;
    mem[11'h39f] = 8'h27;
    mem[11'h3a0] = 8'h30;
    mem[11'h3a1] = 8'h17;
    mem[11'h3a2] = 8'h1b;
    mem[11'h3a3] = 8'h18;
    mem[11'h3a4] = 8'h69;
    mem[11'h3a5] = 8'h27;
    mem[11'h3a6] = 8'h30;
    mem[11'h3a7] = 8'h17;
    mem[11'h3a8] = 8'h1c;
    mem[11'h3a9] = 8'h17;
    mem[11'h3aa] = 8'h69;
    mem[11'h3ab] = 8'h27;
    mem[11'h3ac] = 8'h2f;
    mem[11'h3ad] = 8'h17;
    mem[11'h3ae] = 8'h1d;
    mem[11'h3af] = 8'h18;
    mem[11'h3b0] = 8'h68;
    mem[11'h3b1] = 8'h27;
    mem[11'h3b2] = 8'h2e;
    mem[11'h3b3] = 8'h18;
    mem[11'h3b4] = 8'h1e;
    mem[11'h3b5] = 8'h17;
    mem[11'h3b6] = 8'h68;
    mem[11'h3b7] = 8'h27;
    mem[11'h3b8] = 8'h2e;
    mem[11'h3b9] = 8'h17;
    mem[11'h3ba] = 8'h1f;
    mem[11'h3bb] = 8'h18;
    mem[11'h3bc] = 8'h67;
    mem[11'h3bd] = 8'h27;
    mem[11'h3be] = 8'h2d;
    mem[11'h3bf] = 8'h18;
    mem[11'h3c0] = 8'h20;
    mem[11'h3c1] = 8'h18;
    mem[11'h3c2] = 8'h66;
    mem[11'h3c3] = 8'h27;
    mem[11'h3c4] = 8'h2d;
    mem[11'h3c5] = 8'h17;
    mem[11'h3c6] = 8'h21;
    mem[11'h3c7] = 8'h18;
    mem[11'h3c8] = 8'h66;
    mem[11'h3c9] = 8'h27;
    mem[11'h3ca] = 8'h2c;
    mem[11'h3cb] = 8'h18;
    mem[11'h3cc] = 8'h22;
    mem[11'h3cd] = 8'h18;
    mem[11'h3ce] = 8'h65;
    mem[11'h3cf] = 8'h27;
    mem[11'h3d0] = 8'h2b;
    mem[11'h3d1] = 8'h18;
    mem[11'h3d2] = 8'h23;
    mem[11'h3d3] = 8'h19;
    mem[11'h3d4] = 8'h64;
    mem[11'h3d5] = 8'h27;
    mem[11'h3d6] = 8'h2a;
    mem[11'h3d7] = 8'h19;
    mem[11'h3d8] = 8'h24;
    mem[11'h3d9] = 8'h18;
    mem[11'h3da] = 8'h64;
    mem[11'h3db] = 8'h27;
    mem[11'h3dc] = 8'h2a;
    mem[11'h3dd] = 8'h18;
    mem[11'h3de] = 8'h25;
    mem[11'h3df] = 8'h19;
    mem[11'h3e0] = 8'h63;
    mem[11'h3e1] = 8'h27;
    mem[11'h3e2] = 8'h29;
    mem[11'h3e3] = 8'h19;
    mem[11'h3e4] = 8'h26;
    mem[11'h3e5] = 8'h19;
    mem[11'h3e6] = 8'h62;
    mem[11'h3e7] = 8'h27;
    mem[11'h3e8] = 8'h28;
    mem[11'h3e9] = 8'h19;
    mem[11'h3ea] = 8'h28;
    mem[11'h3eb] = 8'h18;
    mem[11'h3ec] = 8'h62;
    mem[11'h3ed] = 8'h27;
    mem[11'h3ee] = 8'h28;
    mem[11'h3ef] = 8'h19;
    mem[11'h3f0] = 8'h28;
    mem[11'h3f1] = 8'h19;
    mem[11'h3f2] = 8'h61;
    mem[11'h3f3] = 8'h27;
    mem[11'h3f4] = 8'h27;
    mem[11'h3f5] = 8'h19;
    mem[11'h3f6] = 8'h2a;
    mem[11'h3f7] = 8'h19;
    mem[11'h3f8] = 8'h60;
    mem[11'h3f9] = 8'h27;
    mem[11'h3fa] = 8'h26;
    mem[11'h3fb] = 8'h19;
    mem[11'h3fc] = 8'h2b;
    mem[11'h3fd] = 8'h1a;
    mem[11'h3fe] = 8'h5f;
    mem[11'h3ff] = 8'h27;
    mem[11'h400] = 8'h25;
    mem[11'h401] = 8'h1a;
    mem[11'h402] = 8'h2c;
    mem[11'h403] = 8'h1a;
    mem[11'h404] = 8'h5e;
    mem[11'h405] = 8'h27;
    mem[11'h406] = 8'h24;
    mem[11'h407] = 8'h1a;
    mem[11'h408] = 8'h2e;
    mem[11'h409] = 8'h19;
    mem[11'h40a] = 8'h5e;
    mem[11'h40b] = 8'h27;
    mem[11'h40c] = 8'h24;
    mem[11'h40d] = 8'h1a;
    mem[11'h40e] = 8'h2e;
    mem[11'h40f] = 8'h1a;
    mem[11'h410] = 8'h5d;
    mem[11'h411] = 8'h27;
    mem[11'h412] = 8'h23;
    mem[11'h413] = 8'h1a;
    mem[11'h414] = 8'h30;
    mem[11'h415] = 8'h1a;
    mem[11'h416] = 8'h5c;
    mem[11'h417] = 8'h27;
    mem[11'h418] = 8'h22;
    mem[11'h419] = 8'h1a;
    mem[11'h41a] = 8'h32;
    mem[11'h41b] = 8'h1a;
    mem[11'h41c] = 8'h5b;
    mem[11'h41d] = 8'h27;
    mem[11'h41e] = 8'h21;
    mem[11'h41f] = 8'h1b;
    mem[11'h420] = 8'h32;
    mem[11'h421] = 8'h1b;
    mem[11'h422] = 8'h5a;
    mem[11'h423] = 8'h27;
    mem[11'h424] = 8'h20;
    mem[11'h425] = 8'h1b;
    mem[11'h426] = 8'h34;
    mem[11'h427] = 8'h1b;
    mem[11'h428] = 8'h59;
    mem[11'h429] = 8'h27;
    mem[11'h42a] = 8'h1f;
    mem[11'h42b] = 8'h1b;
    mem[11'h42c] = 8'h36;
    mem[11'h42d] = 8'h1b;
    mem[11'h42e] = 8'h58;
    mem[11'h42f] = 8'h27;
    mem[11'h430] = 8'h1e;
    mem[11'h431] = 8'h1b;
    mem[11'h432] = 8'h37;
    mem[11'h433] = 8'h1c;
    mem[11'h434] = 8'h57;
    mem[11'h435] = 8'h27;
    mem[11'h436] = 8'h1d;
    mem[11'h437] = 8'h1c;
    mem[11'h438] = 8'h38;
    mem[11'h439] = 8'h1c;
    mem[11'h43a] = 8'h56;
    mem[11'h43b] = 8'h27;
    mem[11'h43c] = 8'h1c;
    mem[11'h43d] = 8'h1c;
    mem[11'h43e] = 8'h3a;
    mem[11'h43f] = 8'h1c;
    mem[11'h440] = 8'h55;
    mem[11'h441] = 8'h27;
    mem[11'h442] = 8'h1b;
    mem[11'h443] = 8'h1c;
    mem[11'h444] = 8'h3c;
    mem[11'h445] = 8'h1c;
    mem[11'h446] = 8'h54;
    mem[11'h447] = 8'h27;
    mem[11'h448] = 8'h1a;
    mem[11'h449] = 8'h1c;
    mem[11'h44a] = 8'h3e;
    mem[11'h44b] = 8'h1c;
    mem[11'h44c] = 8'h53;
    mem[11'h44d] = 8'h27;
    mem[11'h44e] = 8'h19;
    mem[11'h44f] = 8'h1d;
    mem[11'h450] = 8'h3e;
    mem[11'h451] = 8'h1d;
    mem[11'h452] = 8'h52;
    mem[11'h453] = 8'h27;
    mem[11'h454] = 8'h18;
    mem[11'h455] = 8'h1d;
    mem[11'h456] = 8'h40;
    mem[11'h457] = 8'h1d;
    mem[11'h458] = 8'h51;
    mem[11'h459] = 8'h27;
    mem[11'h45a] = 8'h17;
    mem[11'h45b] = 8'h1d;
    mem[11'h45c] = 8'h42;
    mem[11'h45d] = 8'h1e;
    mem[11'h45e] = 8'h4f;
    mem[11'h45f] = 8'h27;
    mem[11'h460] = 8'h15;
    mem[11'h461] = 8'h1e;
    mem[11'h462] = 8'h44;
    mem[11'h463] = 8'h1e;
    mem[11'h464] = 8'h4e;
    mem[11'h465] = 8'h27;
    mem[11'h466] = 8'h14;
    mem[11'h467] = 8'h1e;
    mem[11'h468] = 8'h46;
    mem[11'h469] = 8'h1e;
    mem[11'h46a] = 8'h4d;
    mem[11'h46b] = 8'h27;
    mem[11'h46c] = 8'h13;
    mem[11'h46d] = 8'h1e;
    mem[11'h46e] = 8'h48;
    mem[11'h46f] = 8'h1e;
    mem[11'h470] = 8'h4c;
    mem[11'h471] = 8'h27;
    mem[11'h472] = 8'h12;
    mem[11'h473] = 8'h1e;
    mem[11'h474] = 8'h49;
    mem[11'h475] = 8'h20;
    mem[11'h476] = 8'h4a;
    mem[11'h477] = 8'h27;
    mem[11'h478] = 8'h10;
    mem[11'h479] = 8'h20;
    mem[11'h47a] = 8'h4a;
    mem[11'h47b] = 8'h20;
    mem[11'h47c] = 8'h49;
    mem[11'h47d] = 8'h27;
    mem[11'h47e] = 8'h0f;
    mem[11'h47f] = 8'h20;
    mem[11'h480] = 8'h4c;
    mem[11'h481] = 8'h21;
    mem[11'h482] = 8'h47;
    mem[11'h483] = 8'h27;
    mem[11'h484] = 8'h0d;
    mem[11'h485] = 8'h21;
    mem[11'h486] = 8'h4e;
    mem[11'h487] = 8'h21;
    mem[11'h488] = 8'h46;
    mem[11'h489] = 8'h27;
    mem[11'h48a] = 8'h0c;
    mem[11'h48b] = 8'h21;
    mem[11'h48c] = 8'h50;
    mem[11'h48d] = 8'h22;
    mem[11'h48e] = 8'h44;
    mem[11'h48f] = 8'h27;
    mem[11'h490] = 8'h0b;
    mem[11'h491] = 8'h21;
    mem[11'h492] = 8'h52;
    mem[11'h493] = 8'h22;
    mem[11'h494] = 8'h43;
    mem[11'h495] = 8'h27;
    mem[11'h496] = 8'h0a;
    mem[11'h497] = 8'h21;
    mem[11'h498] = 8'h54;
    mem[11'h499] = 8'h23;
    mem[11'h49a] = 8'h41;
    mem[11'h49b] = 8'h27;
    mem[11'h49c] = 8'h0a;
    mem[11'h49d] = 8'h20;
    mem[11'h49e] = 8'h56;
    mem[11'h49f] = 8'h24;
    mem[11'h4a0] = 8'h3f;
    mem[11'h4a1] = 8'h27;
    mem[11'h4a2] = 8'h0a;
    mem[11'h4a3] = 8'h1f;
    mem[11'h4a4] = 8'h58;
    mem[11'h4a5] = 8'h24;
    mem[11'h4a6] = 8'h3e;
    mem[11'h4a7] = 8'h27;
    mem[11'h4a8] = 8'h0a;
    mem[11'h4a9] = 8'h1e;
    mem[11'h4aa] = 8'h5b;
    mem[11'h4ab] = 8'h24;
    mem[11'h4ac] = 8'h3c;
    mem[11'h4ad] = 8'h27;
    mem[11'h4ae] = 8'h0a;
    mem[11'h4af] = 8'h1d;
    mem[11'h4b0] = 8'h5d;
    mem[11'h4b1] = 8'h25;
    mem[11'h4b2] = 8'h3a;
    mem[11'h4b3] = 8'h27;
    mem[11'h4b4] = 8'h0a;
    mem[11'h4b5] = 8'h1b;
    mem[11'h4b6] = 8'h60;
    mem[11'h4b7] = 8'h26;
    mem[11'h4b8] = 8'h38;
    mem[11'h4b9] = 8'h27;
    mem[11'h4ba] = 8'h0a;
    mem[11'h4bb] = 8'h1a;
    mem[11'h4bc] = 8'h62;
    mem[11'h4bd] = 8'h27;
    mem[11'h4be] = 8'h36;
    mem[11'h4bf] = 8'h27;
    mem[11'h4c0] = 8'h0a;
    mem[11'h4c1] = 8'h19;
    mem[11'h4c2] = 8'h64;
    mem[11'h4c3] = 8'h29;
    mem[11'h4c4] = 8'h33;
    mem[11'h4c5] = 8'h27;
    mem[11'h4c6] = 8'h0a;
    mem[11'h4c7] = 8'h18;
    mem[11'h4c8] = 8'h67;
    mem[11'h4c9] = 8'h29;
    mem[11'h4ca] = 8'h31;
    mem[11'h4cb] = 8'h27;
    mem[11'h4cc] = 8'h0a;
    mem[11'h4cd] = 8'h17;
    mem[11'h4ce] = 8'h69;
    mem[11'h4cf] = 8'h2b;
    mem[11'h4d0] = 8'h2e;
    mem[11'h4d1] = 8'h27;
    mem[11'h4d2] = 8'h0a;
    mem[11'h4d3] = 8'h15;
    mem[11'h4d4] = 8'h6c;
    mem[11'h4d5] = 8'h2d;
    mem[11'h4d6] = 8'h2b;
    mem[11'h4d7] = 8'h27;
    mem[11'h4d8] = 8'h0a;
    mem[11'h4d9] = 8'h14;
    mem[11'h4da] = 8'h6e;
    mem[11'h4db] = 8'h2f;
    mem[11'h4dc] = 8'h28;
    mem[11'h4dd] = 8'h27;
    mem[11'h4de] = 8'h0a;
    mem[11'h4df] = 8'h13;
    mem[11'h4e0] = 8'h71;
    mem[11'h4e1] = 8'h30;
    mem[11'h4e2] = 8'h25;
    mem[11'h4e3] = 8'h27;
    mem[11'h4e4] = 8'h0a;
    mem[11'h4e5] = 8'h11;
    mem[11'h4e6] = 8'h74;
    mem[11'h4e7] = 8'h33;
    mem[11'h4e8] = 8'h21;
    mem[11'h4e9] = 8'h27;
    mem[11'h4ea] = 8'h0a;
    mem[11'h4eb] = 8'h10;
    mem[11'h4ec] = 8'h77;
    mem[11'h4ed] = 8'h36;
    mem[11'h4ee] = 8'h1c;
    mem[11'h4ef] = 8'h27;
    mem[11'h4f0] = 8'h0a;
    mem[11'h4f1] = 8'h0f;
    mem[11'h4f2] = 8'h79;
    mem[11'h4f3] = 8'h3c;
    mem[11'h4f4] = 8'h15;
    mem[11'h4f5] = 8'h27;
    mem[11'h4f6] = 8'h0a;
    mem[11'h4f7] = 8'h0d;
    mem[11'h4f8] = 8'h7d;
    mem[11'h4f9] = 8'h78;
    mem[11'h4fa] = 8'h0a;
    mem[11'h4fb] = 8'h0c;
    mem[11'h4fc] = 8'h7f;
    mem[11'h4fd] = 8'h77;
    mem[11'h4fe] = 8'h0a;
    mem[11'h4ff] = 8'h0a;
    mem[11'h500] = 8'h83;
    mem[11'h501] = 8'h75;
    mem[11'h502] = 8'h0a;
    mem[11'h503] = 8'h08;
    mem[11'h504] = 8'h87;
    mem[11'h505] = 8'h73;
    mem[11'h506] = 8'h0a;
    mem[11'h507] = 8'h07;
    mem[11'h508] = 8'h89;
    mem[11'h509] = 8'h72;
    mem[11'h50a] = 8'h0a;
    mem[11'h50b] = 8'h05;
    mem[11'h50c] = 8'h8d;
    mem[11'h50d] = 8'h70;
    mem[11'h50e] = 8'h0a;
    mem[11'h50f] = 8'h03;
    mem[11'h510] = 8'h91;
    mem[11'h511] = 8'h6e;
    mem[11'h512] = 8'h0a;
    mem[11'h513] = 8'h01;
    mem[11'h514] = 8'h95;
    mem[11'h515] = 8'h6c;
    mem[11'h516] = 8'ha4;
    mem[11'h517] = 8'h6a;
    mem[11'h518] = 8'ha6;
    mem[11'h519] = 8'h68;
    mem[11'h51a] = 8'ha8;
    mem[11'h51b] = 8'h66;
    mem[11'h51c] = 8'hab;
    mem[11'h51d] = 8'h63;
    mem[11'h51e] = 8'had;
    mem[11'h51f] = 8'h61;
    mem[11'h520] = 8'hb0;
    mem[11'h521] = 8'h5b;
    mem[11'h522] = 8'hb6;
    mem[11'h523] = 8'h55;
    mem[11'h524] = 8'hbc;
    mem[11'h525] = 8'h4f;
    mem[11'h526] = 8'hc2;
    mem[11'h527] = 8'h49;
    mem[11'h528] = 8'hc9;
    mem[11'h529] = 8'h41;
    mem[11'h52a] = 8'hd1;
    mem[11'h52b] = 8'h39;
    mem[11'h52c] = 8'hda;
    mem[11'h52d] = 8'h2f;
    mem[11'h52e] = 8'he5;
    mem[11'h52f] = 8'h22;
    mem[11'h530] = 8'hf9;
    mem[11'h531] = 8'h0a;
  end
  assign len = mem[addr];
endmodule
