
/*
 * Copyright (c) 2024 Tiny Tapeout LTD
 * SPDX-License-Identifier: Apache-2.0
 * Author: Renaldas Zioma
 */

`default_nettype none

// parameter LOGO_SIZE = 272;  // Size of the logo in pixels
parameter LOGO_SIZE = 266;  // Size of the logo in pixels
parameter DISPLAY_WIDTH = 640;  // VGA display width
parameter DISPLAY_HEIGHT = 480;  // VGA display height

// `define ROM1 1

module tt_um_rejunity_vga_logo (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // VGA signals
  wire hsync;
  wire vsync;
  reg [1:0] R;
  reg [1:0] G;
  reg [1:0] B;
  wire video_active;
  wire [9:0] pix_x;
  wire [9:0] pix_y;


  // TinyVGA PMOD
  assign uo_out  = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

  // Unused outputs assigned to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in[7:1], uio_in};

  hvsync_generator vga_sync_gen (
      .clk(clk),
      .reset(~rst_n),
      .hsync(hsync),
      .vsync(vsync),
      .display_on(video_active),
      .hpos(pix_x),
      .vpos(pix_y)
  );

`ifdef ROM1
  wire pixel_value;
  bitmap_rom rom1 (
      .x(pix_x[6:0]),
      .y(pix_y[6:0]),
      .pixel(pixel_value)
  );

  assign {R, G, B } = (video_active&pixel_value) ? 6'b11_11_00 : 6'b00_00_00;

`else
  reg [11:0] addr;
  reg [7:0] len;
  bitmap_rom_rle rom2 (
    .addr(addr),
    .len(len)
  );

  assign {R, G, B } = (video_active&pixel_value&(pix_x<=(LOGO_SIZE))) ? 6'b11_11_00 : 6'b00_00_00;

  // increase couner every frame (vsync happens once per frame)
  reg [7:0] counter;
  reg pixel_value;
  always @(posedge clk) begin
    if (~rst_n) begin
      counter <= 0;
    end else begin
      if (vsync) begin
        addr <= 0;
        counter <= 0;
        pixel_value <= 0;
      end else if (pix_x < LOGO_SIZE && pix_y < LOGO_SIZE) begin
        if (counter >= len) begin
          addr <= addr + 1;
          counter <= 0;
          pixel_value <= ~pixel_value;
        end else begin
          counter <= counter + 1;
        end
      end
    end
  end  
`endif

endmodule

// --------------------------------------------------------

module bitmap_rom (
    input wire [6:0] x,
    input wire [6:0] y,
    output wire pixel
);

  reg [7:0] mem[2047:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h80;
    mem[23] = 8'hff;
    mem[24] = 8'hff;
    mem[25] = 8'h01;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'hfc;
    mem[39] = 8'hff;
    mem[40] = 8'hff;
    mem[41] = 8'h3f;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'hc0;
    mem[54] = 8'hff;
    mem[55] = 8'hff;
    mem[56] = 8'hff;
    mem[57] = 8'hff;
    mem[58] = 8'h03;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'hf8;
    mem[70] = 8'hff;
    mem[71] = 8'hff;
    mem[72] = 8'hff;
    mem[73] = 8'hff;
    mem[74] = 8'h1f;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'hff;
    mem[86] = 8'hff;
    mem[87] = 8'hff;
    mem[88] = 8'hff;
    mem[89] = 8'hff;
    mem[90] = 8'hff;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'hc0;
    mem[101] = 8'hff;
    mem[102] = 8'hff;
    mem[103] = 8'hff;
    mem[104] = 8'hff;
    mem[105] = 8'hff;
    mem[106] = 8'hff;
    mem[107] = 8'h03;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'hf0;
    mem[117] = 8'hff;
    mem[118] = 8'hff;
    mem[119] = 8'hff;
    mem[120] = 8'hff;
    mem[121] = 8'hff;
    mem[122] = 8'hff;
    mem[123] = 8'h0f;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'hfc;
    mem[133] = 8'hff;
    mem[134] = 8'hff;
    mem[135] = 8'hff;
    mem[136] = 8'hff;
    mem[137] = 8'hff;
    mem[138] = 8'hff;
    mem[139] = 8'h3f;
    mem[140] = 8'h00;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'hff;
    mem[149] = 8'hff;
    mem[150] = 8'hff;
    mem[151] = 8'hff;
    mem[152] = 8'hff;
    mem[153] = 8'hff;
    mem[154] = 8'hff;
    mem[155] = 8'hff;
    mem[156] = 8'h00;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h00;
    mem[162] = 8'h00;
    mem[163] = 8'hc0;
    mem[164] = 8'hff;
    mem[165] = 8'hff;
    mem[166] = 8'hff;
    mem[167] = 8'hff;
    mem[168] = 8'hff;
    mem[169] = 8'hff;
    mem[170] = 8'hff;
    mem[171] = 8'hff;
    mem[172] = 8'h03;
    mem[173] = 8'h00;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h00;
    mem[178] = 8'h00;
    mem[179] = 8'he0;
    mem[180] = 8'hff;
    mem[181] = 8'hff;
    mem[182] = 8'hff;
    mem[183] = 8'h7f;
    mem[184] = 8'hfe;
    mem[185] = 8'hff;
    mem[186] = 8'hff;
    mem[187] = 8'hff;
    mem[188] = 8'h07;
    mem[189] = 8'h00;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
    mem[192] = 8'h00;
    mem[193] = 8'h00;
    mem[194] = 8'h00;
    mem[195] = 8'hf8;
    mem[196] = 8'hff;
    mem[197] = 8'hff;
    mem[198] = 8'h3f;
    mem[199] = 8'h00;
    mem[200] = 8'h00;
    mem[201] = 8'hfc;
    mem[202] = 8'hff;
    mem[203] = 8'hff;
    mem[204] = 8'h1f;
    mem[205] = 8'h00;
    mem[206] = 8'h00;
    mem[207] = 8'h00;
    mem[208] = 8'h00;
    mem[209] = 8'h00;
    mem[210] = 8'h00;
    mem[211] = 8'hfc;
    mem[212] = 8'hff;
    mem[213] = 8'hff;
    mem[214] = 8'h03;
    mem[215] = 8'h00;
    mem[216] = 8'h00;
    mem[217] = 8'hc0;
    mem[218] = 8'hff;
    mem[219] = 8'hff;
    mem[220] = 8'h3f;
    mem[221] = 8'h00;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'h00;
    mem[227] = 8'hfe;
    mem[228] = 8'hff;
    mem[229] = 8'h7f;
    mem[230] = 8'h00;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'hfe;
    mem[235] = 8'hff;
    mem[236] = 8'h7f;
    mem[237] = 8'h00;
    mem[238] = 8'h00;
    mem[239] = 8'h00;
    mem[240] = 8'h00;
    mem[241] = 8'h00;
    mem[242] = 8'h80;
    mem[243] = 8'hff;
    mem[244] = 8'hff;
    mem[245] = 8'h0f;
    mem[246] = 8'h00;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'hf0;
    mem[251] = 8'hff;
    mem[252] = 8'hff;
    mem[253] = 8'h01;
    mem[254] = 8'h00;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'h00;
    mem[258] = 8'hc0;
    mem[259] = 8'hff;
    mem[260] = 8'hff;
    mem[261] = 8'h03;
    mem[262] = 8'h00;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'hc0;
    mem[267] = 8'hff;
    mem[268] = 8'hff;
    mem[269] = 8'h03;
    mem[270] = 8'h00;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'he0;
    mem[275] = 8'hff;
    mem[276] = 8'hff;
    mem[277] = 8'h00;
    mem[278] = 8'h00;
    mem[279] = 8'h00;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'h00;
    mem[283] = 8'hff;
    mem[284] = 8'hff;
    mem[285] = 8'h07;
    mem[286] = 8'h00;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'hf0;
    mem[291] = 8'hff;
    mem[292] = 8'h3f;
    mem[293] = 8'h00;
    mem[294] = 8'h00;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'h00;
    mem[299] = 8'hfc;
    mem[300] = 8'hff;
    mem[301] = 8'h0f;
    mem[302] = 8'h00;
    mem[303] = 8'h00;
    mem[304] = 8'h00;
    mem[305] = 8'h00;
    mem[306] = 8'hf8;
    mem[307] = 8'hff;
    mem[308] = 8'h0f;
    mem[309] = 8'h00;
    mem[310] = 8'h00;
    mem[311] = 8'h00;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'h00;
    mem[315] = 8'hf0;
    mem[316] = 8'hff;
    mem[317] = 8'h1f;
    mem[318] = 8'h00;
    mem[319] = 8'h00;
    mem[320] = 8'h00;
    mem[321] = 8'h00;
    mem[322] = 8'hfc;
    mem[323] = 8'hff;
    mem[324] = 8'h07;
    mem[325] = 8'h00;
    mem[326] = 8'h00;
    mem[327] = 8'h00;
    mem[328] = 8'h00;
    mem[329] = 8'h00;
    mem[330] = 8'h00;
    mem[331] = 8'he0;
    mem[332] = 8'hff;
    mem[333] = 8'h3f;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
    mem[336] = 8'h00;
    mem[337] = 8'h00;
    mem[338] = 8'hfe;
    mem[339] = 8'hff;
    mem[340] = 8'h01;
    mem[341] = 8'h00;
    mem[342] = 8'h00;
    mem[343] = 8'h00;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'h00;
    mem[347] = 8'h80;
    mem[348] = 8'hff;
    mem[349] = 8'h7f;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'h00;
    mem[354] = 8'hff;
    mem[355] = 8'hff;
    mem[356] = 8'h00;
    mem[357] = 8'h00;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'hff;
    mem[365] = 8'hff;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h80;
    mem[370] = 8'hff;
    mem[371] = 8'h7f;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'hfe;
    mem[381] = 8'hff;
    mem[382] = 8'h01;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h80;
    mem[386] = 8'hff;
    mem[387] = 8'h3f;
    mem[388] = 8'h00;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'hfc;
    mem[397] = 8'hff;
    mem[398] = 8'h01;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'hc0;
    mem[402] = 8'hff;
    mem[403] = 8'h1f;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'hf8;
    mem[413] = 8'hff;
    mem[414] = 8'h03;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'he0;
    mem[418] = 8'hff;
    mem[419] = 8'h0f;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'he0;
    mem[429] = 8'hff;
    mem[430] = 8'h07;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'hf0;
    mem[434] = 8'hff;
    mem[435] = 8'hff;
    mem[436] = 8'hff;
    mem[437] = 8'hff;
    mem[438] = 8'hff;
    mem[439] = 8'hff;
    mem[440] = 8'hff;
    mem[441] = 8'h0f;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'hc0;
    mem[445] = 8'hff;
    mem[446] = 8'h0f;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'hf0;
    mem[450] = 8'hff;
    mem[451] = 8'hff;
    mem[452] = 8'hff;
    mem[453] = 8'hff;
    mem[454] = 8'hff;
    mem[455] = 8'hff;
    mem[456] = 8'hff;
    mem[457] = 8'h0f;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'hc0;
    mem[461] = 8'hff;
    mem[462] = 8'h0f;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'hf8;
    mem[466] = 8'hff;
    mem[467] = 8'hff;
    mem[468] = 8'hff;
    mem[469] = 8'hff;
    mem[470] = 8'hff;
    mem[471] = 8'hff;
    mem[472] = 8'hff;
    mem[473] = 8'h0f;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h80;
    mem[477] = 8'hff;
    mem[478] = 8'h1f;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'hfc;
    mem[482] = 8'hff;
    mem[483] = 8'hff;
    mem[484] = 8'hff;
    mem[485] = 8'hff;
    mem[486] = 8'hff;
    mem[487] = 8'hff;
    mem[488] = 8'hff;
    mem[489] = 8'h0f;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'hff;
    mem[494] = 8'h3f;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'hfc;
    mem[498] = 8'hff;
    mem[499] = 8'hff;
    mem[500] = 8'hff;
    mem[501] = 8'hff;
    mem[502] = 8'hff;
    mem[503] = 8'hff;
    mem[504] = 8'hff;
    mem[505] = 8'h0f;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'hfe;
    mem[510] = 8'h3f;
    mem[511] = 8'h00;
    mem[512] = 8'h00;
    mem[513] = 8'hfe;
    mem[514] = 8'hff;
    mem[515] = 8'hff;
    mem[516] = 8'hff;
    mem[517] = 8'hff;
    mem[518] = 8'hff;
    mem[519] = 8'hff;
    mem[520] = 8'hff;
    mem[521] = 8'h0f;
    mem[522] = 8'h00;
    mem[523] = 8'h00;
    mem[524] = 8'h00;
    mem[525] = 8'hfc;
    mem[526] = 8'h7f;
    mem[527] = 8'h00;
    mem[528] = 8'h00;
    mem[529] = 8'hfe;
    mem[530] = 8'hff;
    mem[531] = 8'hff;
    mem[532] = 8'hff;
    mem[533] = 8'hff;
    mem[534] = 8'hff;
    mem[535] = 8'hff;
    mem[536] = 8'hff;
    mem[537] = 8'h0f;
    mem[538] = 8'h00;
    mem[539] = 8'h00;
    mem[540] = 8'h00;
    mem[541] = 8'hf8;
    mem[542] = 8'h7f;
    mem[543] = 8'h00;
    mem[544] = 8'h00;
    mem[545] = 8'hff;
    mem[546] = 8'hff;
    mem[547] = 8'hff;
    mem[548] = 8'hff;
    mem[549] = 8'hff;
    mem[550] = 8'hff;
    mem[551] = 8'hff;
    mem[552] = 8'hff;
    mem[553] = 8'h0f;
    mem[554] = 8'h00;
    mem[555] = 8'h00;
    mem[556] = 8'h00;
    mem[557] = 8'hf8;
    mem[558] = 8'hff;
    mem[559] = 8'h00;
    mem[560] = 8'h00;
    mem[561] = 8'hff;
    mem[562] = 8'hff;
    mem[563] = 8'hff;
    mem[564] = 8'hff;
    mem[565] = 8'hff;
    mem[566] = 8'hff;
    mem[567] = 8'hff;
    mem[568] = 8'hff;
    mem[569] = 8'h0f;
    mem[570] = 8'h00;
    mem[571] = 8'h00;
    mem[572] = 8'h00;
    mem[573] = 8'hf0;
    mem[574] = 8'hff;
    mem[575] = 8'h00;
    mem[576] = 8'h80;
    mem[577] = 8'hff;
    mem[578] = 8'hff;
    mem[579] = 8'hff;
    mem[580] = 8'hff;
    mem[581] = 8'hff;
    mem[582] = 8'hff;
    mem[583] = 8'hff;
    mem[584] = 8'hff;
    mem[585] = 8'h0f;
    mem[586] = 8'h00;
    mem[587] = 8'h00;
    mem[588] = 8'h00;
    mem[589] = 8'he0;
    mem[590] = 8'hff;
    mem[591] = 8'h01;
    mem[592] = 8'h80;
    mem[593] = 8'hff;
    mem[594] = 8'hff;
    mem[595] = 8'hff;
    mem[596] = 8'hff;
    mem[597] = 8'hff;
    mem[598] = 8'hff;
    mem[599] = 8'hff;
    mem[600] = 8'hff;
    mem[601] = 8'h0f;
    mem[602] = 8'h00;
    mem[603] = 8'h00;
    mem[604] = 8'h00;
    mem[605] = 8'he0;
    mem[606] = 8'hff;
    mem[607] = 8'h01;
    mem[608] = 8'hc0;
    mem[609] = 8'hff;
    mem[610] = 8'hff;
    mem[611] = 8'hff;
    mem[612] = 8'hff;
    mem[613] = 8'hff;
    mem[614] = 8'hff;
    mem[615] = 8'hff;
    mem[616] = 8'hff;
    mem[617] = 8'h0f;
    mem[618] = 8'h00;
    mem[619] = 8'h00;
    mem[620] = 8'h00;
    mem[621] = 8'hc0;
    mem[622] = 8'hff;
    mem[623] = 8'h03;
    mem[624] = 8'hc0;
    mem[625] = 8'hff;
    mem[626] = 8'hff;
    mem[627] = 8'hff;
    mem[628] = 8'hff;
    mem[629] = 8'hff;
    mem[630] = 8'hff;
    mem[631] = 8'hff;
    mem[632] = 8'hff;
    mem[633] = 8'h0f;
    mem[634] = 8'h00;
    mem[635] = 8'h00;
    mem[636] = 8'h00;
    mem[637] = 8'hc0;
    mem[638] = 8'hff;
    mem[639] = 8'h03;
    mem[640] = 8'he0;
    mem[641] = 8'hff;
    mem[642] = 8'hff;
    mem[643] = 8'hff;
    mem[644] = 8'hff;
    mem[645] = 8'hff;
    mem[646] = 8'hff;
    mem[647] = 8'hff;
    mem[648] = 8'hff;
    mem[649] = 8'h0f;
    mem[650] = 8'h00;
    mem[651] = 8'h00;
    mem[652] = 8'h00;
    mem[653] = 8'h80;
    mem[654] = 8'hff;
    mem[655] = 8'h07;
    mem[656] = 8'he0;
    mem[657] = 8'hff;
    mem[658] = 8'hff;
    mem[659] = 8'hff;
    mem[660] = 8'hff;
    mem[661] = 8'hff;
    mem[662] = 8'hff;
    mem[663] = 8'hff;
    mem[664] = 8'hff;
    mem[665] = 8'h0f;
    mem[666] = 8'h00;
    mem[667] = 8'h00;
    mem[668] = 8'h00;
    mem[669] = 8'h80;
    mem[670] = 8'hff;
    mem[671] = 8'h07;
    mem[672] = 8'he0;
    mem[673] = 8'hff;
    mem[674] = 8'hff;
    mem[675] = 8'hff;
    mem[676] = 8'hff;
    mem[677] = 8'hff;
    mem[678] = 8'hff;
    mem[679] = 8'hff;
    mem[680] = 8'hff;
    mem[681] = 8'h0f;
    mem[682] = 8'h00;
    mem[683] = 8'h00;
    mem[684] = 8'h00;
    mem[685] = 8'h00;
    mem[686] = 8'hff;
    mem[687] = 8'h07;
    mem[688] = 8'hf0;
    mem[689] = 8'hff;
    mem[690] = 8'hff;
    mem[691] = 8'hff;
    mem[692] = 8'hff;
    mem[693] = 8'hff;
    mem[694] = 8'hff;
    mem[695] = 8'hff;
    mem[696] = 8'hff;
    mem[697] = 8'h0f;
    mem[698] = 8'h00;
    mem[699] = 8'h00;
    mem[700] = 8'h00;
    mem[701] = 8'h00;
    mem[702] = 8'hff;
    mem[703] = 8'h0f;
    mem[704] = 8'hf0;
    mem[705] = 8'hff;
    mem[706] = 8'hff;
    mem[707] = 8'hff;
    mem[708] = 8'hff;
    mem[709] = 8'hff;
    mem[710] = 8'hff;
    mem[711] = 8'hff;
    mem[712] = 8'hff;
    mem[713] = 8'h0f;
    mem[714] = 8'h00;
    mem[715] = 8'h00;
    mem[716] = 8'h00;
    mem[717] = 8'h00;
    mem[718] = 8'hfe;
    mem[719] = 8'h0f;
    mem[720] = 8'h00;
    mem[721] = 8'h00;
    mem[722] = 8'h00;
    mem[723] = 8'h00;
    mem[724] = 8'h80;
    mem[725] = 8'hff;
    mem[726] = 8'hff;
    mem[727] = 8'h03;
    mem[728] = 8'h00;
    mem[729] = 8'h00;
    mem[730] = 8'h00;
    mem[731] = 8'h00;
    mem[732] = 8'h00;
    mem[733] = 8'h00;
    mem[734] = 8'hfe;
    mem[735] = 8'h0f;
    mem[736] = 8'h00;
    mem[737] = 8'h00;
    mem[738] = 8'h00;
    mem[739] = 8'h00;
    mem[740] = 8'h80;
    mem[741] = 8'hff;
    mem[742] = 8'hff;
    mem[743] = 8'h03;
    mem[744] = 8'h00;
    mem[745] = 8'h00;
    mem[746] = 8'h00;
    mem[747] = 8'h00;
    mem[748] = 8'h00;
    mem[749] = 8'h00;
    mem[750] = 8'hfe;
    mem[751] = 8'h1f;
    mem[752] = 8'h00;
    mem[753] = 8'h00;
    mem[754] = 8'h00;
    mem[755] = 8'h00;
    mem[756] = 8'h80;
    mem[757] = 8'hff;
    mem[758] = 8'hff;
    mem[759] = 8'h03;
    mem[760] = 8'h00;
    mem[761] = 8'h00;
    mem[762] = 8'h00;
    mem[763] = 8'h00;
    mem[764] = 8'h00;
    mem[765] = 8'h00;
    mem[766] = 8'hfc;
    mem[767] = 8'h1f;
    mem[768] = 8'h00;
    mem[769] = 8'h00;
    mem[770] = 8'h00;
    mem[771] = 8'h00;
    mem[772] = 8'h80;
    mem[773] = 8'hff;
    mem[774] = 8'hff;
    mem[775] = 8'h03;
    mem[776] = 8'h00;
    mem[777] = 8'h00;
    mem[778] = 8'h00;
    mem[779] = 8'h00;
    mem[780] = 8'h00;
    mem[781] = 8'h00;
    mem[782] = 8'hfc;
    mem[783] = 8'h1f;
    mem[784] = 8'h00;
    mem[785] = 8'h00;
    mem[786] = 8'h00;
    mem[787] = 8'h00;
    mem[788] = 8'h80;
    mem[789] = 8'hff;
    mem[790] = 8'hff;
    mem[791] = 8'h03;
    mem[792] = 8'h00;
    mem[793] = 8'h00;
    mem[794] = 8'h00;
    mem[795] = 8'h00;
    mem[796] = 8'h00;
    mem[797] = 8'h00;
    mem[798] = 8'hfc;
    mem[799] = 8'h3f;
    mem[800] = 8'hfc;
    mem[801] = 8'h1f;
    mem[802] = 8'h00;
    mem[803] = 8'h00;
    mem[804] = 8'h80;
    mem[805] = 8'hff;
    mem[806] = 8'hff;
    mem[807] = 8'h03;
    mem[808] = 8'h00;
    mem[809] = 8'h00;
    mem[810] = 8'h00;
    mem[811] = 8'h00;
    mem[812] = 8'h00;
    mem[813] = 8'h00;
    mem[814] = 8'hf8;
    mem[815] = 8'h3f;
    mem[816] = 8'hfc;
    mem[817] = 8'h1f;
    mem[818] = 8'h00;
    mem[819] = 8'h00;
    mem[820] = 8'h80;
    mem[821] = 8'hff;
    mem[822] = 8'hff;
    mem[823] = 8'h03;
    mem[824] = 8'h00;
    mem[825] = 8'h00;
    mem[826] = 8'h00;
    mem[827] = 8'h00;
    mem[828] = 8'h00;
    mem[829] = 8'h00;
    mem[830] = 8'hf8;
    mem[831] = 8'h3f;
    mem[832] = 8'hfc;
    mem[833] = 8'h1f;
    mem[834] = 8'h00;
    mem[835] = 8'h00;
    mem[836] = 8'h80;
    mem[837] = 8'hff;
    mem[838] = 8'hff;
    mem[839] = 8'h03;
    mem[840] = 8'h00;
    mem[841] = 8'h00;
    mem[842] = 8'h00;
    mem[843] = 8'h00;
    mem[844] = 8'h00;
    mem[845] = 8'h00;
    mem[846] = 8'hf8;
    mem[847] = 8'h3f;
    mem[848] = 8'hfc;
    mem[849] = 8'h1f;
    mem[850] = 8'h00;
    mem[851] = 8'h00;
    mem[852] = 8'h80;
    mem[853] = 8'hff;
    mem[854] = 8'hff;
    mem[855] = 8'h03;
    mem[856] = 8'h00;
    mem[857] = 8'h00;
    mem[858] = 8'h00;
    mem[859] = 8'h00;
    mem[860] = 8'h00;
    mem[861] = 8'h00;
    mem[862] = 8'hf8;
    mem[863] = 8'h3f;
    mem[864] = 8'hfc;
    mem[865] = 8'h0f;
    mem[866] = 8'h00;
    mem[867] = 8'h00;
    mem[868] = 8'h80;
    mem[869] = 8'hff;
    mem[870] = 8'hff;
    mem[871] = 8'h03;
    mem[872] = 8'h00;
    mem[873] = 8'h00;
    mem[874] = 8'h00;
    mem[875] = 8'h00;
    mem[876] = 8'h00;
    mem[877] = 8'h00;
    mem[878] = 8'hf0;
    mem[879] = 8'h3f;
    mem[880] = 8'hfe;
    mem[881] = 8'h0f;
    mem[882] = 8'h00;
    mem[883] = 8'h00;
    mem[884] = 8'h80;
    mem[885] = 8'hff;
    mem[886] = 8'hff;
    mem[887] = 8'h03;
    mem[888] = 8'h00;
    mem[889] = 8'h00;
    mem[890] = 8'h00;
    mem[891] = 8'h00;
    mem[892] = 8'h00;
    mem[893] = 8'h00;
    mem[894] = 8'hf0;
    mem[895] = 8'h7f;
    mem[896] = 8'hfe;
    mem[897] = 8'h0f;
    mem[898] = 8'h00;
    mem[899] = 8'h00;
    mem[900] = 8'h80;
    mem[901] = 8'hff;
    mem[902] = 8'hff;
    mem[903] = 8'h03;
    mem[904] = 8'h00;
    mem[905] = 8'h00;
    mem[906] = 8'h00;
    mem[907] = 8'h00;
    mem[908] = 8'h00;
    mem[909] = 8'h00;
    mem[910] = 8'hf0;
    mem[911] = 8'h7f;
    mem[912] = 8'hfe;
    mem[913] = 8'h0f;
    mem[914] = 8'h00;
    mem[915] = 8'h00;
    mem[916] = 8'h80;
    mem[917] = 8'hff;
    mem[918] = 8'hff;
    mem[919] = 8'h03;
    mem[920] = 8'h00;
    mem[921] = 8'h00;
    mem[922] = 8'h00;
    mem[923] = 8'h00;
    mem[924] = 8'h00;
    mem[925] = 8'h00;
    mem[926] = 8'hf0;
    mem[927] = 8'h7f;
    mem[928] = 8'hfe;
    mem[929] = 8'h0f;
    mem[930] = 8'h00;
    mem[931] = 8'h00;
    mem[932] = 8'h80;
    mem[933] = 8'hff;
    mem[934] = 8'hff;
    mem[935] = 8'hff;
    mem[936] = 8'hff;
    mem[937] = 8'hff;
    mem[938] = 8'hff;
    mem[939] = 8'hff;
    mem[940] = 8'hff;
    mem[941] = 8'h01;
    mem[942] = 8'hf0;
    mem[943] = 8'h7f;
    mem[944] = 8'hfe;
    mem[945] = 8'h0f;
    mem[946] = 8'h00;
    mem[947] = 8'h00;
    mem[948] = 8'h80;
    mem[949] = 8'hff;
    mem[950] = 8'hff;
    mem[951] = 8'hff;
    mem[952] = 8'hff;
    mem[953] = 8'hff;
    mem[954] = 8'hff;
    mem[955] = 8'hff;
    mem[956] = 8'hff;
    mem[957] = 8'h01;
    mem[958] = 8'hf0;
    mem[959] = 8'h7f;
    mem[960] = 8'hfe;
    mem[961] = 8'h0f;
    mem[962] = 8'h00;
    mem[963] = 8'h00;
    mem[964] = 8'h80;
    mem[965] = 8'hff;
    mem[966] = 8'hff;
    mem[967] = 8'hff;
    mem[968] = 8'hff;
    mem[969] = 8'hff;
    mem[970] = 8'hff;
    mem[971] = 8'hff;
    mem[972] = 8'hff;
    mem[973] = 8'h01;
    mem[974] = 8'hf0;
    mem[975] = 8'h7f;
    mem[976] = 8'hfe;
    mem[977] = 8'h07;
    mem[978] = 8'h00;
    mem[979] = 8'h00;
    mem[980] = 8'h80;
    mem[981] = 8'hff;
    mem[982] = 8'hff;
    mem[983] = 8'hff;
    mem[984] = 8'hff;
    mem[985] = 8'hff;
    mem[986] = 8'hff;
    mem[987] = 8'hff;
    mem[988] = 8'hff;
    mem[989] = 8'h01;
    mem[990] = 8'hf0;
    mem[991] = 8'h7f;
    mem[992] = 8'hfe;
    mem[993] = 8'h07;
    mem[994] = 8'h00;
    mem[995] = 8'h00;
    mem[996] = 8'h80;
    mem[997] = 8'hff;
    mem[998] = 8'hff;
    mem[999] = 8'hff;
    mem[1000] = 8'hff;
    mem[1001] = 8'hff;
    mem[1002] = 8'hff;
    mem[1003] = 8'hff;
    mem[1004] = 8'hff;
    mem[1005] = 8'h01;
    mem[1006] = 8'hf0;
    mem[1007] = 8'h7f;
    mem[1008] = 8'hfe;
    mem[1009] = 8'h07;
    mem[1010] = 8'h00;
    mem[1011] = 8'h00;
    mem[1012] = 8'h80;
    mem[1013] = 8'hff;
    mem[1014] = 8'hff;
    mem[1015] = 8'hff;
    mem[1016] = 8'hff;
    mem[1017] = 8'hff;
    mem[1018] = 8'hff;
    mem[1019] = 8'hff;
    mem[1020] = 8'hff;
    mem[1021] = 8'h01;
    mem[1022] = 8'he0;
    mem[1023] = 8'h7f;
    mem[1024] = 8'hfe;
    mem[1025] = 8'h07;
    mem[1026] = 8'h00;
    mem[1027] = 8'h00;
    mem[1028] = 8'h80;
    mem[1029] = 8'hff;
    mem[1030] = 8'hff;
    mem[1031] = 8'hff;
    mem[1032] = 8'hff;
    mem[1033] = 8'hff;
    mem[1034] = 8'hff;
    mem[1035] = 8'hff;
    mem[1036] = 8'hff;
    mem[1037] = 8'h01;
    mem[1038] = 8'he0;
    mem[1039] = 8'h7f;
    mem[1040] = 8'hfe;
    mem[1041] = 8'h07;
    mem[1042] = 8'h00;
    mem[1043] = 8'h00;
    mem[1044] = 8'h80;
    mem[1045] = 8'hff;
    mem[1046] = 8'hff;
    mem[1047] = 8'hff;
    mem[1048] = 8'hff;
    mem[1049] = 8'hff;
    mem[1050] = 8'hff;
    mem[1051] = 8'hff;
    mem[1052] = 8'hff;
    mem[1053] = 8'h01;
    mem[1054] = 8'he0;
    mem[1055] = 8'h7f;
    mem[1056] = 8'hfe;
    mem[1057] = 8'h0f;
    mem[1058] = 8'h00;
    mem[1059] = 8'h00;
    mem[1060] = 8'h80;
    mem[1061] = 8'hff;
    mem[1062] = 8'hff;
    mem[1063] = 8'hff;
    mem[1064] = 8'hff;
    mem[1065] = 8'hff;
    mem[1066] = 8'hff;
    mem[1067] = 8'hff;
    mem[1068] = 8'hff;
    mem[1069] = 8'h01;
    mem[1070] = 8'hf0;
    mem[1071] = 8'h7f;
    mem[1072] = 8'hfe;
    mem[1073] = 8'h0f;
    mem[1074] = 8'h00;
    mem[1075] = 8'h00;
    mem[1076] = 8'h80;
    mem[1077] = 8'hff;
    mem[1078] = 8'hff;
    mem[1079] = 8'hff;
    mem[1080] = 8'hff;
    mem[1081] = 8'hff;
    mem[1082] = 8'hff;
    mem[1083] = 8'hff;
    mem[1084] = 8'hff;
    mem[1085] = 8'h01;
    mem[1086] = 8'hf0;
    mem[1087] = 8'h7f;
    mem[1088] = 8'hfe;
    mem[1089] = 8'h0f;
    mem[1090] = 8'h00;
    mem[1091] = 8'h00;
    mem[1092] = 8'h80;
    mem[1093] = 8'hff;
    mem[1094] = 8'hff;
    mem[1095] = 8'hff;
    mem[1096] = 8'hff;
    mem[1097] = 8'hff;
    mem[1098] = 8'hff;
    mem[1099] = 8'hff;
    mem[1100] = 8'hff;
    mem[1101] = 8'h01;
    mem[1102] = 8'hf0;
    mem[1103] = 8'h7f;
    mem[1104] = 8'hfe;
    mem[1105] = 8'h0f;
    mem[1106] = 8'h00;
    mem[1107] = 8'h00;
    mem[1108] = 8'h80;
    mem[1109] = 8'hff;
    mem[1110] = 8'hff;
    mem[1111] = 8'hff;
    mem[1112] = 8'hff;
    mem[1113] = 8'hff;
    mem[1114] = 8'hff;
    mem[1115] = 8'hff;
    mem[1116] = 8'hff;
    mem[1117] = 8'h01;
    mem[1118] = 8'hf0;
    mem[1119] = 8'h7f;
    mem[1120] = 8'hfe;
    mem[1121] = 8'h0f;
    mem[1122] = 8'h00;
    mem[1123] = 8'h00;
    mem[1124] = 8'h80;
    mem[1125] = 8'hff;
    mem[1126] = 8'hff;
    mem[1127] = 8'hff;
    mem[1128] = 8'hff;
    mem[1129] = 8'hff;
    mem[1130] = 8'hff;
    mem[1131] = 8'hff;
    mem[1132] = 8'hff;
    mem[1133] = 8'h01;
    mem[1134] = 8'hf0;
    mem[1135] = 8'h7f;
    mem[1136] = 8'hfe;
    mem[1137] = 8'h0f;
    mem[1138] = 8'h00;
    mem[1139] = 8'h00;
    mem[1140] = 8'h80;
    mem[1141] = 8'hff;
    mem[1142] = 8'hff;
    mem[1143] = 8'hff;
    mem[1144] = 8'hff;
    mem[1145] = 8'hff;
    mem[1146] = 8'hff;
    mem[1147] = 8'hff;
    mem[1148] = 8'hff;
    mem[1149] = 8'h01;
    mem[1150] = 8'hf0;
    mem[1151] = 8'h7f;
    mem[1152] = 8'hfe;
    mem[1153] = 8'h0f;
    mem[1154] = 8'h00;
    mem[1155] = 8'h00;
    mem[1156] = 8'h80;
    mem[1157] = 8'hff;
    mem[1158] = 8'hff;
    mem[1159] = 8'hff;
    mem[1160] = 8'hff;
    mem[1161] = 8'hff;
    mem[1162] = 8'hff;
    mem[1163] = 8'hff;
    mem[1164] = 8'hff;
    mem[1165] = 8'h01;
    mem[1166] = 8'hf0;
    mem[1167] = 8'h7f;
    mem[1168] = 8'hfc;
    mem[1169] = 8'h0f;
    mem[1170] = 8'h00;
    mem[1171] = 8'h00;
    mem[1172] = 8'h80;
    mem[1173] = 8'hff;
    mem[1174] = 8'hff;
    mem[1175] = 8'hff;
    mem[1176] = 8'hff;
    mem[1177] = 8'hff;
    mem[1178] = 8'hff;
    mem[1179] = 8'hff;
    mem[1180] = 8'hff;
    mem[1181] = 8'h01;
    mem[1182] = 8'hf0;
    mem[1183] = 8'h3f;
    mem[1184] = 8'hfc;
    mem[1185] = 8'h1f;
    mem[1186] = 8'h00;
    mem[1187] = 8'h00;
    mem[1188] = 8'h80;
    mem[1189] = 8'hff;
    mem[1190] = 8'hff;
    mem[1191] = 8'hff;
    mem[1192] = 8'hff;
    mem[1193] = 8'hff;
    mem[1194] = 8'hff;
    mem[1195] = 8'hff;
    mem[1196] = 8'hff;
    mem[1197] = 8'h01;
    mem[1198] = 8'hf8;
    mem[1199] = 8'h3f;
    mem[1200] = 8'hfc;
    mem[1201] = 8'h1f;
    mem[1202] = 8'h00;
    mem[1203] = 8'h00;
    mem[1204] = 8'h80;
    mem[1205] = 8'hff;
    mem[1206] = 8'hff;
    mem[1207] = 8'hff;
    mem[1208] = 8'hff;
    mem[1209] = 8'hff;
    mem[1210] = 8'hff;
    mem[1211] = 8'hff;
    mem[1212] = 8'hff;
    mem[1213] = 8'h01;
    mem[1214] = 8'hf8;
    mem[1215] = 8'h3f;
    mem[1216] = 8'hfc;
    mem[1217] = 8'h1f;
    mem[1218] = 8'h00;
    mem[1219] = 8'h00;
    mem[1220] = 8'h80;
    mem[1221] = 8'hff;
    mem[1222] = 8'hff;
    mem[1223] = 8'h03;
    mem[1224] = 8'hf0;
    mem[1225] = 8'hff;
    mem[1226] = 8'h7f;
    mem[1227] = 8'h00;
    mem[1228] = 8'h00;
    mem[1229] = 8'h00;
    mem[1230] = 8'hf8;
    mem[1231] = 8'h3f;
    mem[1232] = 8'hfc;
    mem[1233] = 8'h1f;
    mem[1234] = 8'h00;
    mem[1235] = 8'h00;
    mem[1236] = 8'h80;
    mem[1237] = 8'hff;
    mem[1238] = 8'hff;
    mem[1239] = 8'h03;
    mem[1240] = 8'hf0;
    mem[1241] = 8'hff;
    mem[1242] = 8'h7f;
    mem[1243] = 8'h00;
    mem[1244] = 8'h00;
    mem[1245] = 8'h00;
    mem[1246] = 8'hf8;
    mem[1247] = 8'h3f;
    mem[1248] = 8'hfc;
    mem[1249] = 8'h3f;
    mem[1250] = 8'h00;
    mem[1251] = 8'h00;
    mem[1252] = 8'h80;
    mem[1253] = 8'hff;
    mem[1254] = 8'hff;
    mem[1255] = 8'h03;
    mem[1256] = 8'hf0;
    mem[1257] = 8'hff;
    mem[1258] = 8'h7f;
    mem[1259] = 8'h00;
    mem[1260] = 8'h00;
    mem[1261] = 8'h00;
    mem[1262] = 8'hfc;
    mem[1263] = 8'h3f;
    mem[1264] = 8'hf8;
    mem[1265] = 8'h3f;
    mem[1266] = 8'h00;
    mem[1267] = 8'h00;
    mem[1268] = 8'h80;
    mem[1269] = 8'hff;
    mem[1270] = 8'hff;
    mem[1271] = 8'h03;
    mem[1272] = 8'hf0;
    mem[1273] = 8'hff;
    mem[1274] = 8'h7f;
    mem[1275] = 8'h00;
    mem[1276] = 8'h00;
    mem[1277] = 8'h00;
    mem[1278] = 8'hfc;
    mem[1279] = 8'h1f;
    mem[1280] = 8'hf8;
    mem[1281] = 8'h3f;
    mem[1282] = 8'h00;
    mem[1283] = 8'h00;
    mem[1284] = 8'h80;
    mem[1285] = 8'hff;
    mem[1286] = 8'hff;
    mem[1287] = 8'h03;
    mem[1288] = 8'hf0;
    mem[1289] = 8'hff;
    mem[1290] = 8'h7f;
    mem[1291] = 8'h00;
    mem[1292] = 8'h00;
    mem[1293] = 8'h00;
    mem[1294] = 8'hfc;
    mem[1295] = 8'h1f;
    mem[1296] = 8'hf8;
    mem[1297] = 8'h7f;
    mem[1298] = 8'h00;
    mem[1299] = 8'h00;
    mem[1300] = 8'h80;
    mem[1301] = 8'hff;
    mem[1302] = 8'hff;
    mem[1303] = 8'h03;
    mem[1304] = 8'hf0;
    mem[1305] = 8'hff;
    mem[1306] = 8'h7f;
    mem[1307] = 8'h00;
    mem[1308] = 8'h00;
    mem[1309] = 8'h00;
    mem[1310] = 8'hfe;
    mem[1311] = 8'h1f;
    mem[1312] = 8'hf0;
    mem[1313] = 8'h7f;
    mem[1314] = 8'h00;
    mem[1315] = 8'h00;
    mem[1316] = 8'h80;
    mem[1317] = 8'hff;
    mem[1318] = 8'hff;
    mem[1319] = 8'h03;
    mem[1320] = 8'hf0;
    mem[1321] = 8'hff;
    mem[1322] = 8'h7f;
    mem[1323] = 8'h00;
    mem[1324] = 8'h00;
    mem[1325] = 8'h00;
    mem[1326] = 8'hfe;
    mem[1327] = 8'h0f;
    mem[1328] = 8'hf0;
    mem[1329] = 8'h7f;
    mem[1330] = 8'h00;
    mem[1331] = 8'h00;
    mem[1332] = 8'h80;
    mem[1333] = 8'hff;
    mem[1334] = 8'hff;
    mem[1335] = 8'h03;
    mem[1336] = 8'hf0;
    mem[1337] = 8'hff;
    mem[1338] = 8'h7f;
    mem[1339] = 8'h00;
    mem[1340] = 8'h00;
    mem[1341] = 8'h00;
    mem[1342] = 8'hfe;
    mem[1343] = 8'h0f;
    mem[1344] = 8'hf0;
    mem[1345] = 8'hff;
    mem[1346] = 8'h00;
    mem[1347] = 8'h00;
    mem[1348] = 8'h80;
    mem[1349] = 8'hff;
    mem[1350] = 8'hff;
    mem[1351] = 8'h03;
    mem[1352] = 8'hf0;
    mem[1353] = 8'hff;
    mem[1354] = 8'h7f;
    mem[1355] = 8'h00;
    mem[1356] = 8'h00;
    mem[1357] = 8'h00;
    mem[1358] = 8'hff;
    mem[1359] = 8'h0f;
    mem[1360] = 8'he0;
    mem[1361] = 8'hff;
    mem[1362] = 8'h00;
    mem[1363] = 8'h00;
    mem[1364] = 8'h80;
    mem[1365] = 8'hff;
    mem[1366] = 8'hff;
    mem[1367] = 8'h03;
    mem[1368] = 8'hf0;
    mem[1369] = 8'hff;
    mem[1370] = 8'h7f;
    mem[1371] = 8'h00;
    mem[1372] = 8'h00;
    mem[1373] = 8'h00;
    mem[1374] = 8'hff;
    mem[1375] = 8'h07;
    mem[1376] = 8'he0;
    mem[1377] = 8'hff;
    mem[1378] = 8'h01;
    mem[1379] = 8'h00;
    mem[1380] = 8'h80;
    mem[1381] = 8'hff;
    mem[1382] = 8'hff;
    mem[1383] = 8'h03;
    mem[1384] = 8'hf0;
    mem[1385] = 8'hff;
    mem[1386] = 8'h7f;
    mem[1387] = 8'h00;
    mem[1388] = 8'h00;
    mem[1389] = 8'h80;
    mem[1390] = 8'hff;
    mem[1391] = 8'h07;
    mem[1392] = 8'he0;
    mem[1393] = 8'hff;
    mem[1394] = 8'h01;
    mem[1395] = 8'h00;
    mem[1396] = 8'h00;
    mem[1397] = 8'h00;
    mem[1398] = 8'h00;
    mem[1399] = 8'h00;
    mem[1400] = 8'hf0;
    mem[1401] = 8'hff;
    mem[1402] = 8'h7f;
    mem[1403] = 8'h00;
    mem[1404] = 8'h00;
    mem[1405] = 8'h80;
    mem[1406] = 8'hff;
    mem[1407] = 8'h07;
    mem[1408] = 8'hc0;
    mem[1409] = 8'hff;
    mem[1410] = 8'h03;
    mem[1411] = 8'h00;
    mem[1412] = 8'h00;
    mem[1413] = 8'h00;
    mem[1414] = 8'h00;
    mem[1415] = 8'h00;
    mem[1416] = 8'hf0;
    mem[1417] = 8'hff;
    mem[1418] = 8'h7f;
    mem[1419] = 8'h00;
    mem[1420] = 8'h00;
    mem[1421] = 8'hc0;
    mem[1422] = 8'hff;
    mem[1423] = 8'h03;
    mem[1424] = 8'hc0;
    mem[1425] = 8'hff;
    mem[1426] = 8'h03;
    mem[1427] = 8'h00;
    mem[1428] = 8'h00;
    mem[1429] = 8'h00;
    mem[1430] = 8'h00;
    mem[1431] = 8'h00;
    mem[1432] = 8'hf0;
    mem[1433] = 8'hff;
    mem[1434] = 8'h7f;
    mem[1435] = 8'h00;
    mem[1436] = 8'h00;
    mem[1437] = 8'hc0;
    mem[1438] = 8'hff;
    mem[1439] = 8'h03;
    mem[1440] = 8'h80;
    mem[1441] = 8'hff;
    mem[1442] = 8'h07;
    mem[1443] = 8'h00;
    mem[1444] = 8'h00;
    mem[1445] = 8'h00;
    mem[1446] = 8'h00;
    mem[1447] = 8'h00;
    mem[1448] = 8'hf0;
    mem[1449] = 8'hff;
    mem[1450] = 8'h7f;
    mem[1451] = 8'h00;
    mem[1452] = 8'h00;
    mem[1453] = 8'he0;
    mem[1454] = 8'hff;
    mem[1455] = 8'h01;
    mem[1456] = 8'h80;
    mem[1457] = 8'hff;
    mem[1458] = 8'h07;
    mem[1459] = 8'h00;
    mem[1460] = 8'h00;
    mem[1461] = 8'h00;
    mem[1462] = 8'h00;
    mem[1463] = 8'h00;
    mem[1464] = 8'hf0;
    mem[1465] = 8'hff;
    mem[1466] = 8'h7f;
    mem[1467] = 8'h00;
    mem[1468] = 8'h00;
    mem[1469] = 8'he0;
    mem[1470] = 8'hff;
    mem[1471] = 8'h01;
    mem[1472] = 8'h00;
    mem[1473] = 8'hff;
    mem[1474] = 8'h0f;
    mem[1475] = 8'h00;
    mem[1476] = 8'h00;
    mem[1477] = 8'h00;
    mem[1478] = 8'h00;
    mem[1479] = 8'h00;
    mem[1480] = 8'hf0;
    mem[1481] = 8'hff;
    mem[1482] = 8'h7f;
    mem[1483] = 8'h00;
    mem[1484] = 8'h00;
    mem[1485] = 8'hf0;
    mem[1486] = 8'hff;
    mem[1487] = 8'h00;
    mem[1488] = 8'h00;
    mem[1489] = 8'hff;
    mem[1490] = 8'h1f;
    mem[1491] = 8'h00;
    mem[1492] = 8'h00;
    mem[1493] = 8'h00;
    mem[1494] = 8'h00;
    mem[1495] = 8'h00;
    mem[1496] = 8'hf0;
    mem[1497] = 8'hff;
    mem[1498] = 8'h7f;
    mem[1499] = 8'h00;
    mem[1500] = 8'h00;
    mem[1501] = 8'hf8;
    mem[1502] = 8'hff;
    mem[1503] = 8'h00;
    mem[1504] = 8'h00;
    mem[1505] = 8'hfe;
    mem[1506] = 8'h1f;
    mem[1507] = 8'h00;
    mem[1508] = 8'h00;
    mem[1509] = 8'h00;
    mem[1510] = 8'h00;
    mem[1511] = 8'h00;
    mem[1512] = 8'hf0;
    mem[1513] = 8'hff;
    mem[1514] = 8'h7f;
    mem[1515] = 8'h00;
    mem[1516] = 8'h00;
    mem[1517] = 8'hf8;
    mem[1518] = 8'h7f;
    mem[1519] = 8'h00;
    mem[1520] = 8'h00;
    mem[1521] = 8'hfe;
    mem[1522] = 8'h3f;
    mem[1523] = 8'h00;
    mem[1524] = 8'h00;
    mem[1525] = 8'h00;
    mem[1526] = 8'h00;
    mem[1527] = 8'h00;
    mem[1528] = 8'hf0;
    mem[1529] = 8'hff;
    mem[1530] = 8'h7f;
    mem[1531] = 8'h00;
    mem[1532] = 8'h00;
    mem[1533] = 8'hfc;
    mem[1534] = 8'h7f;
    mem[1535] = 8'h00;
    mem[1536] = 8'h00;
    mem[1537] = 8'hfc;
    mem[1538] = 8'h7f;
    mem[1539] = 8'h00;
    mem[1540] = 8'h00;
    mem[1541] = 8'h00;
    mem[1542] = 8'h00;
    mem[1543] = 8'h00;
    mem[1544] = 8'hf0;
    mem[1545] = 8'hff;
    mem[1546] = 8'h7f;
    mem[1547] = 8'h00;
    mem[1548] = 8'h00;
    mem[1549] = 8'hfe;
    mem[1550] = 8'h3f;
    mem[1551] = 8'h00;
    mem[1552] = 8'h00;
    mem[1553] = 8'hfc;
    mem[1554] = 8'hff;
    mem[1555] = 8'h00;
    mem[1556] = 8'h00;
    mem[1557] = 8'h00;
    mem[1558] = 8'h00;
    mem[1559] = 8'h00;
    mem[1560] = 8'hf0;
    mem[1561] = 8'hff;
    mem[1562] = 8'h7f;
    mem[1563] = 8'h00;
    mem[1564] = 8'h00;
    mem[1565] = 8'hff;
    mem[1566] = 8'h3f;
    mem[1567] = 8'h00;
    mem[1568] = 8'h00;
    mem[1569] = 8'hf8;
    mem[1570] = 8'hff;
    mem[1571] = 8'h01;
    mem[1572] = 8'h00;
    mem[1573] = 8'h00;
    mem[1574] = 8'h00;
    mem[1575] = 8'h00;
    mem[1576] = 8'hf0;
    mem[1577] = 8'hff;
    mem[1578] = 8'h7f;
    mem[1579] = 8'h00;
    mem[1580] = 8'h80;
    mem[1581] = 8'hff;
    mem[1582] = 8'h1f;
    mem[1583] = 8'h00;
    mem[1584] = 8'h00;
    mem[1585] = 8'hf0;
    mem[1586] = 8'hff;
    mem[1587] = 8'h03;
    mem[1588] = 8'h00;
    mem[1589] = 8'h00;
    mem[1590] = 8'h00;
    mem[1591] = 8'h00;
    mem[1592] = 8'hf0;
    mem[1593] = 8'hff;
    mem[1594] = 8'h7f;
    mem[1595] = 8'h00;
    mem[1596] = 8'hc0;
    mem[1597] = 8'hff;
    mem[1598] = 8'h0f;
    mem[1599] = 8'h00;
    mem[1600] = 8'h00;
    mem[1601] = 8'hf0;
    mem[1602] = 8'hff;
    mem[1603] = 8'h03;
    mem[1604] = 8'h00;
    mem[1605] = 8'h00;
    mem[1606] = 8'h00;
    mem[1607] = 8'h00;
    mem[1608] = 8'hf0;
    mem[1609] = 8'hff;
    mem[1610] = 8'h7f;
    mem[1611] = 8'h00;
    mem[1612] = 8'hc0;
    mem[1613] = 8'hff;
    mem[1614] = 8'h0f;
    mem[1615] = 8'h00;
    mem[1616] = 8'h00;
    mem[1617] = 8'he0;
    mem[1618] = 8'hff;
    mem[1619] = 8'h07;
    mem[1620] = 8'h00;
    mem[1621] = 8'h00;
    mem[1622] = 8'h00;
    mem[1623] = 8'h00;
    mem[1624] = 8'hf0;
    mem[1625] = 8'hff;
    mem[1626] = 8'h7f;
    mem[1627] = 8'h00;
    mem[1628] = 8'he0;
    mem[1629] = 8'hff;
    mem[1630] = 8'h07;
    mem[1631] = 8'h00;
    mem[1632] = 8'h00;
    mem[1633] = 8'hc0;
    mem[1634] = 8'hff;
    mem[1635] = 8'h1f;
    mem[1636] = 8'h00;
    mem[1637] = 8'h00;
    mem[1638] = 8'h00;
    mem[1639] = 8'h00;
    mem[1640] = 8'hf0;
    mem[1641] = 8'hff;
    mem[1642] = 8'h7f;
    mem[1643] = 8'h00;
    mem[1644] = 8'hf0;
    mem[1645] = 8'hff;
    mem[1646] = 8'h03;
    mem[1647] = 8'h00;
    mem[1648] = 8'h00;
    mem[1649] = 8'h80;
    mem[1650] = 8'hff;
    mem[1651] = 8'h3f;
    mem[1652] = 8'h00;
    mem[1653] = 8'h00;
    mem[1654] = 8'h00;
    mem[1655] = 8'h00;
    mem[1656] = 8'hf0;
    mem[1657] = 8'hff;
    mem[1658] = 8'h7f;
    mem[1659] = 8'h00;
    mem[1660] = 8'hfc;
    mem[1661] = 8'hff;
    mem[1662] = 8'h01;
    mem[1663] = 8'h00;
    mem[1664] = 8'h00;
    mem[1665] = 8'h80;
    mem[1666] = 8'hff;
    mem[1667] = 8'h7f;
    mem[1668] = 8'h00;
    mem[1669] = 8'h00;
    mem[1670] = 8'h00;
    mem[1671] = 8'h00;
    mem[1672] = 8'hf0;
    mem[1673] = 8'hff;
    mem[1674] = 8'h7f;
    mem[1675] = 8'h00;
    mem[1676] = 8'hfe;
    mem[1677] = 8'hff;
    mem[1678] = 8'h01;
    mem[1679] = 8'h00;
    mem[1680] = 8'h00;
    mem[1681] = 8'h00;
    mem[1682] = 8'hff;
    mem[1683] = 8'hff;
    mem[1684] = 8'h00;
    mem[1685] = 8'h00;
    mem[1686] = 8'h00;
    mem[1687] = 8'h00;
    mem[1688] = 8'hf0;
    mem[1689] = 8'hff;
    mem[1690] = 8'h7f;
    mem[1691] = 8'h00;
    mem[1692] = 8'hff;
    mem[1693] = 8'hff;
    mem[1694] = 8'h00;
    mem[1695] = 8'h00;
    mem[1696] = 8'h00;
    mem[1697] = 8'h00;
    mem[1698] = 8'hfe;
    mem[1699] = 8'hff;
    mem[1700] = 8'h01;
    mem[1701] = 8'h00;
    mem[1702] = 8'h00;
    mem[1703] = 8'h00;
    mem[1704] = 8'hf0;
    mem[1705] = 8'hff;
    mem[1706] = 8'h7f;
    mem[1707] = 8'h80;
    mem[1708] = 8'hff;
    mem[1709] = 8'h7f;
    mem[1710] = 8'h00;
    mem[1711] = 8'h00;
    mem[1712] = 8'h00;
    mem[1713] = 8'h00;
    mem[1714] = 8'hfc;
    mem[1715] = 8'hff;
    mem[1716] = 8'h07;
    mem[1717] = 8'h00;
    mem[1718] = 8'h00;
    mem[1719] = 8'h00;
    mem[1720] = 8'hf0;
    mem[1721] = 8'hff;
    mem[1722] = 8'h7f;
    mem[1723] = 8'he0;
    mem[1724] = 8'hff;
    mem[1725] = 8'h3f;
    mem[1726] = 8'h00;
    mem[1727] = 8'h00;
    mem[1728] = 8'h00;
    mem[1729] = 8'h00;
    mem[1730] = 8'hf8;
    mem[1731] = 8'hff;
    mem[1732] = 8'h0f;
    mem[1733] = 8'h00;
    mem[1734] = 8'h00;
    mem[1735] = 8'h00;
    mem[1736] = 8'hf0;
    mem[1737] = 8'hff;
    mem[1738] = 8'h7f;
    mem[1739] = 8'hf0;
    mem[1740] = 8'hff;
    mem[1741] = 8'h1f;
    mem[1742] = 8'h00;
    mem[1743] = 8'h00;
    mem[1744] = 8'h00;
    mem[1745] = 8'h00;
    mem[1746] = 8'hf0;
    mem[1747] = 8'hff;
    mem[1748] = 8'h3f;
    mem[1749] = 8'h00;
    mem[1750] = 8'h00;
    mem[1751] = 8'h00;
    mem[1752] = 8'hf0;
    mem[1753] = 8'hff;
    mem[1754] = 8'h7f;
    mem[1755] = 8'hf0;
    mem[1756] = 8'hff;
    mem[1757] = 8'h0f;
    mem[1758] = 8'h00;
    mem[1759] = 8'h00;
    mem[1760] = 8'h00;
    mem[1761] = 8'h00;
    mem[1762] = 8'he0;
    mem[1763] = 8'hff;
    mem[1764] = 8'hff;
    mem[1765] = 8'h00;
    mem[1766] = 8'h00;
    mem[1767] = 8'h00;
    mem[1768] = 8'hf0;
    mem[1769] = 8'hff;
    mem[1770] = 8'h7f;
    mem[1771] = 8'hf0;
    mem[1772] = 8'hff;
    mem[1773] = 8'h07;
    mem[1774] = 8'h00;
    mem[1775] = 8'h00;
    mem[1776] = 8'h00;
    mem[1777] = 8'h00;
    mem[1778] = 8'hc0;
    mem[1779] = 8'hff;
    mem[1780] = 8'hff;
    mem[1781] = 8'h03;
    mem[1782] = 8'h00;
    mem[1783] = 8'h00;
    mem[1784] = 8'hf0;
    mem[1785] = 8'hff;
    mem[1786] = 8'h7f;
    mem[1787] = 8'hf0;
    mem[1788] = 8'hff;
    mem[1789] = 8'h03;
    mem[1790] = 8'h00;
    mem[1791] = 8'h00;
    mem[1792] = 8'h00;
    mem[1793] = 8'h00;
    mem[1794] = 8'h80;
    mem[1795] = 8'hff;
    mem[1796] = 8'hff;
    mem[1797] = 8'h0f;
    mem[1798] = 8'h00;
    mem[1799] = 8'h00;
    mem[1800] = 8'hf0;
    mem[1801] = 8'hff;
    mem[1802] = 8'h7f;
    mem[1803] = 8'hf0;
    mem[1804] = 8'hff;
    mem[1805] = 8'h01;
    mem[1806] = 8'h00;
    mem[1807] = 8'h00;
    mem[1808] = 8'h00;
    mem[1809] = 8'h00;
    mem[1810] = 8'h00;
    mem[1811] = 8'hfe;
    mem[1812] = 8'hff;
    mem[1813] = 8'h7f;
    mem[1814] = 8'h00;
    mem[1815] = 8'h00;
    mem[1816] = 8'hf0;
    mem[1817] = 8'hff;
    mem[1818] = 8'h7f;
    mem[1819] = 8'hf0;
    mem[1820] = 8'h7f;
    mem[1821] = 8'h00;
    mem[1822] = 8'h00;
    mem[1823] = 8'h00;
    mem[1824] = 8'h00;
    mem[1825] = 8'h00;
    mem[1826] = 8'h00;
    mem[1827] = 8'hfc;
    mem[1828] = 8'hff;
    mem[1829] = 8'hff;
    mem[1830] = 8'h03;
    mem[1831] = 8'h00;
    mem[1832] = 8'hf0;
    mem[1833] = 8'hff;
    mem[1834] = 8'h7f;
    mem[1835] = 8'hf0;
    mem[1836] = 8'h3f;
    mem[1837] = 8'h00;
    mem[1838] = 8'h00;
    mem[1839] = 8'h00;
    mem[1840] = 8'h00;
    mem[1841] = 8'h00;
    mem[1842] = 8'h00;
    mem[1843] = 8'hf8;
    mem[1844] = 8'hff;
    mem[1845] = 8'hff;
    mem[1846] = 8'h3f;
    mem[1847] = 8'h00;
    mem[1848] = 8'hf0;
    mem[1849] = 8'hff;
    mem[1850] = 8'h7f;
    mem[1851] = 8'hf0;
    mem[1852] = 8'h1f;
    mem[1853] = 8'h00;
    mem[1854] = 8'h00;
    mem[1855] = 8'h00;
    mem[1856] = 8'h00;
    mem[1857] = 8'h00;
    mem[1858] = 8'h00;
    mem[1859] = 8'he0;
    mem[1860] = 8'hff;
    mem[1861] = 8'hff;
    mem[1862] = 8'hff;
    mem[1863] = 8'h7f;
    mem[1864] = 8'hfc;
    mem[1865] = 8'hff;
    mem[1866] = 8'h7f;
    mem[1867] = 8'hf0;
    mem[1868] = 8'h07;
    mem[1869] = 8'h00;
    mem[1870] = 8'h00;
    mem[1871] = 8'h00;
    mem[1872] = 8'h00;
    mem[1873] = 8'h00;
    mem[1874] = 8'h00;
    mem[1875] = 8'hc0;
    mem[1876] = 8'hff;
    mem[1877] = 8'hff;
    mem[1878] = 8'hff;
    mem[1879] = 8'hff;
    mem[1880] = 8'hff;
    mem[1881] = 8'hff;
    mem[1882] = 8'h7f;
    mem[1883] = 8'hf0;
    mem[1884] = 8'h03;
    mem[1885] = 8'h00;
    mem[1886] = 8'h00;
    mem[1887] = 8'h00;
    mem[1888] = 8'h00;
    mem[1889] = 8'h00;
    mem[1890] = 8'h00;
    mem[1891] = 8'h00;
    mem[1892] = 8'hff;
    mem[1893] = 8'hff;
    mem[1894] = 8'hff;
    mem[1895] = 8'hff;
    mem[1896] = 8'hff;
    mem[1897] = 8'hff;
    mem[1898] = 8'h7f;
    mem[1899] = 8'hf0;
    mem[1900] = 8'h00;
    mem[1901] = 8'h00;
    mem[1902] = 8'h00;
    mem[1903] = 8'h00;
    mem[1904] = 8'h00;
    mem[1905] = 8'h00;
    mem[1906] = 8'h00;
    mem[1907] = 8'h00;
    mem[1908] = 8'hfc;
    mem[1909] = 8'hff;
    mem[1910] = 8'hff;
    mem[1911] = 8'hff;
    mem[1912] = 8'hff;
    mem[1913] = 8'hff;
    mem[1914] = 8'h7f;
    mem[1915] = 8'h30;
    mem[1916] = 8'h00;
    mem[1917] = 8'h00;
    mem[1918] = 8'h00;
    mem[1919] = 8'h00;
    mem[1920] = 8'h00;
    mem[1921] = 8'h00;
    mem[1922] = 8'h00;
    mem[1923] = 8'h00;
    mem[1924] = 8'hf0;
    mem[1925] = 8'hff;
    mem[1926] = 8'hff;
    mem[1927] = 8'hff;
    mem[1928] = 8'hff;
    mem[1929] = 8'hff;
    mem[1930] = 8'h7f;
    mem[1931] = 8'h00;
    mem[1932] = 8'h00;
    mem[1933] = 8'h00;
    mem[1934] = 8'h00;
    mem[1935] = 8'h00;
    mem[1936] = 8'h00;
    mem[1937] = 8'h00;
    mem[1938] = 8'h00;
    mem[1939] = 8'h00;
    mem[1940] = 8'hc0;
    mem[1941] = 8'hff;
    mem[1942] = 8'hff;
    mem[1943] = 8'hff;
    mem[1944] = 8'hff;
    mem[1945] = 8'hff;
    mem[1946] = 8'h7f;
    mem[1947] = 8'h00;
    mem[1948] = 8'h00;
    mem[1949] = 8'h00;
    mem[1950] = 8'h00;
    mem[1951] = 8'h00;
    mem[1952] = 8'h00;
    mem[1953] = 8'h00;
    mem[1954] = 8'h00;
    mem[1955] = 8'h00;
    mem[1956] = 8'h00;
    mem[1957] = 8'hff;
    mem[1958] = 8'hff;
    mem[1959] = 8'hff;
    mem[1960] = 8'hff;
    mem[1961] = 8'hff;
    mem[1962] = 8'h7f;
    mem[1963] = 8'h00;
    mem[1964] = 8'h00;
    mem[1965] = 8'h00;
    mem[1966] = 8'h00;
    mem[1967] = 8'h00;
    mem[1968] = 8'h00;
    mem[1969] = 8'h00;
    mem[1970] = 8'h00;
    mem[1971] = 8'h00;
    mem[1972] = 8'h00;
    mem[1973] = 8'hf8;
    mem[1974] = 8'hff;
    mem[1975] = 8'hff;
    mem[1976] = 8'hff;
    mem[1977] = 8'hff;
    mem[1978] = 8'h1f;
    mem[1979] = 8'h00;
    mem[1980] = 8'h00;
    mem[1981] = 8'h00;
    mem[1982] = 8'h00;
    mem[1983] = 8'h00;
    mem[1984] = 8'h00;
    mem[1985] = 8'h00;
    mem[1986] = 8'h00;
    mem[1987] = 8'h00;
    mem[1988] = 8'h00;
    mem[1989] = 8'hc0;
    mem[1990] = 8'hff;
    mem[1991] = 8'hff;
    mem[1992] = 8'hff;
    mem[1993] = 8'hff;
    mem[1994] = 8'h03;
    mem[1995] = 8'h00;
    mem[1996] = 8'h00;
    mem[1997] = 8'h00;
    mem[1998] = 8'h00;
    mem[1999] = 8'h00;
    mem[2000] = 8'h00;
    mem[2001] = 8'h00;
    mem[2002] = 8'h00;
    mem[2003] = 8'h00;
    mem[2004] = 8'h00;
    mem[2005] = 8'h00;
    mem[2006] = 8'hfc;
    mem[2007] = 8'hff;
    mem[2008] = 8'hff;
    mem[2009] = 8'h3f;
    mem[2010] = 8'h00;
    mem[2011] = 8'h00;
    mem[2012] = 8'h00;
    mem[2013] = 8'h00;
    mem[2014] = 8'h00;
    mem[2015] = 8'h00;
    mem[2016] = 8'h00;
    mem[2017] = 8'h00;
    mem[2018] = 8'h00;
    mem[2019] = 8'h00;
    mem[2020] = 8'h00;
    mem[2021] = 8'h00;
    mem[2022] = 8'h80;
    mem[2023] = 8'hff;
    mem[2024] = 8'hff;
    mem[2025] = 8'h01;
    mem[2026] = 8'h00;
    mem[2027] = 8'h00;
    mem[2028] = 8'h00;
    mem[2029] = 8'h00;
    mem[2030] = 8'h00;
    mem[2031] = 8'h00;
    mem[2032] = 8'h00;
    mem[2033] = 8'h00;
    mem[2034] = 8'h00;
    mem[2035] = 8'h00;
    mem[2036] = 8'h00;
    mem[2037] = 8'h00;
    mem[2038] = 8'h00;
    mem[2039] = 8'h00;
    mem[2040] = 8'h00;
    mem[2041] = 8'h00;
    mem[2042] = 8'h00;
    mem[2043] = 8'h00;
    mem[2044] = 8'h00;
    mem[2045] = 8'h00;
    mem[2046] = 8'h00;
    mem[2047] = 8'h00;
  end

  wire [10:0] addr = {y[6:0], x[6:3]};
  assign pixel = mem[addr][x&7];

endmodule

module bitmap_rom_rle (
    input wire [11:0] addr,
    output wire [7:0] len
);

  reg [7:0] mem[1258:0];
  initial begin
    mem[11'h000] = 8'h73;
    mem[11'h001] = 8'h23;
    mem[11'h002] = 8'hdf;
    mem[11'h003] = 8'h2f;
    mem[11'h004] = 8'hd4;
    mem[11'h005] = 8'h39;
    mem[11'h006] = 8'hcb;
    mem[11'h007] = 8'h41;
    mem[11'h008] = 8'hc3;
    mem[11'h009] = 8'h49;
    mem[11'h00a] = 8'hbc;
    mem[11'h00b] = 8'h4f;
    mem[11'h00c] = 8'hb6;
    mem[11'h00d] = 8'h55;
    mem[11'h00e] = 8'hb0;
    mem[11'h00f] = 8'h5b;
    mem[11'h010] = 8'haa;
    mem[11'h011] = 8'h61;
    mem[11'h012] = 8'ha5;
    mem[11'h013] = 8'h65;
    mem[11'h014] = 8'ha0;
    mem[11'h015] = 8'h6b;
    mem[11'h016] = 8'h9b;
    mem[11'h017] = 8'h6f;
    mem[11'h018] = 8'h97;
    mem[11'h019] = 8'h73;
    mem[11'h01a] = 8'h93;
    mem[11'h01b] = 8'h77;
    mem[11'h01c] = 8'h8f;
    mem[11'h01d] = 8'h7b;
    mem[11'h01e] = 8'h8b;
    mem[11'h01f] = 8'h7f;
    mem[11'h020] = 8'h87;
    mem[11'h021] = 8'h83;
    mem[11'h022] = 8'h84;
    mem[11'h023] = 8'h85;
    mem[11'h024] = 8'h81;
    mem[11'h025] = 8'h89;
    mem[11'h026] = 8'h7d;
    mem[11'h027] = 8'h8d;
    mem[11'h028] = 8'h7a;
    mem[11'h029] = 8'h8f;
    mem[11'h02a] = 8'h77;
    mem[11'h02b] = 8'h3c;
    mem[11'h02c] = 8'h1a;
    mem[11'h02d] = 8'h3b;
    mem[11'h02e] = 8'h74;
    mem[11'h02f] = 8'h36;
    mem[11'h030] = 8'h27;
    mem[11'h031] = 8'h36;
    mem[11'h032] = 8'h71;
    mem[11'h033] = 8'h33;
    mem[11'h034] = 8'h31;
    mem[11'h035] = 8'h33;
    mem[11'h036] = 8'h6e;
    mem[11'h037] = 8'h30;
    mem[11'h038] = 8'h39;
    mem[11'h039] = 8'h30;
    mem[11'h03a] = 8'h6c;
    mem[11'h03b] = 8'h2e;
    mem[11'h03c] = 8'h3f;
    mem[11'h03d] = 8'h2f;
    mem[11'h03e] = 8'h68;
    mem[11'h03f] = 8'h2d;
    mem[11'h040] = 8'h46;
    mem[11'h041] = 8'h2c;
    mem[11'h042] = 8'h66;
    mem[11'h043] = 8'h2b;
    mem[11'h044] = 8'h4b;
    mem[11'h045] = 8'h2b;
    mem[11'h046] = 8'h64;
    mem[11'h047] = 8'h29;
    mem[11'h048] = 8'h51;
    mem[11'h049] = 8'h29;
    mem[11'h04a] = 8'h61;
    mem[11'h04b] = 8'h29;
    mem[11'h04c] = 8'h56;
    mem[11'h04d] = 8'h28;
    mem[11'h04e] = 8'h5e;
    mem[11'h04f] = 8'h27;
    mem[11'h050] = 8'h5b;
    mem[11'h051] = 8'h27;
    mem[11'h052] = 8'h5c;
    mem[11'h053] = 8'h26;
    mem[11'h054] = 8'h5f;
    mem[11'h055] = 8'h26;
    mem[11'h056] = 8'h5a;
    mem[11'h057] = 8'h25;
    mem[11'h058] = 8'h63;
    mem[11'h059] = 8'h25;
    mem[11'h05a] = 8'h58;
    mem[11'h05b] = 8'h24;
    mem[11'h05c] = 8'h67;
    mem[11'h05d] = 8'h24;
    mem[11'h05e] = 8'h56;
    mem[11'h05f] = 8'h23;
    mem[11'h060] = 8'h6b;
    mem[11'h061] = 8'h24;
    mem[11'h062] = 8'h53;
    mem[11'h063] = 8'h23;
    mem[11'h064] = 8'h6e;
    mem[11'h065] = 8'h23;
    mem[11'h066] = 8'h51;
    mem[11'h067] = 8'h22;
    mem[11'h068] = 8'h71;
    mem[11'h069] = 8'h23;
    mem[11'h06a] = 8'h4e;
    mem[11'h06b] = 8'h22;
    mem[11'h06c] = 8'h75;
    mem[11'h06d] = 8'h22;
    mem[11'h06e] = 8'h4c;
    mem[11'h06f] = 8'h22;
    mem[11'h070] = 8'h77;
    mem[11'h071] = 8'h22;
    mem[11'h072] = 8'h4b;
    mem[11'h073] = 8'h20;
    mem[11'h074] = 8'h7b;
    mem[11'h075] = 8'h21;
    mem[11'h076] = 8'h49;
    mem[11'h077] = 8'h20;
    mem[11'h078] = 8'h7d;
    mem[11'h079] = 8'h21;
    mem[11'h07a] = 8'h47;
    mem[11'h07b] = 8'h1f;
    mem[11'h07c] = 8'h81;
    mem[11'h07d] = 8'h20;
    mem[11'h07e] = 8'h45;
    mem[11'h07f] = 8'h1f;
    mem[11'h080] = 8'h83;
    mem[11'h081] = 8'h20;
    mem[11'h082] = 8'h43;
    mem[11'h083] = 8'h1e;
    mem[11'h084] = 8'h87;
    mem[11'h085] = 8'h1e;
    mem[11'h086] = 8'h42;
    mem[11'h087] = 8'h1e;
    mem[11'h088] = 8'h89;
    mem[11'h089] = 8'h1e;
    mem[11'h08a] = 8'h40;
    mem[11'h08b] = 8'h1e;
    mem[11'h08c] = 8'h8b;
    mem[11'h08d] = 8'h1e;
    mem[11'h08e] = 8'h3e;
    mem[11'h08f] = 8'h1e;
    mem[11'h090] = 8'h8d;
    mem[11'h091] = 8'h1e;
    mem[11'h092] = 8'h3c;
    mem[11'h093] = 8'h1d;
    mem[11'h094] = 8'h91;
    mem[11'h095] = 8'h1d;
    mem[11'h096] = 8'h3a;
    mem[11'h097] = 8'h1d;
    mem[11'h098] = 8'h93;
    mem[11'h099] = 8'h1d;
    mem[11'h09a] = 8'h39;
    mem[11'h09b] = 8'h1c;
    mem[11'h09c] = 8'h95;
    mem[11'h09d] = 8'h1c;
    mem[11'h09e] = 8'h38;
    mem[11'h09f] = 8'h1c;
    mem[11'h0a0] = 8'h97;
    mem[11'h0a1] = 8'h1c;
    mem[11'h0a2] = 8'h36;
    mem[11'h0a3] = 8'h1c;
    mem[11'h0a4] = 8'h99;
    mem[11'h0a5] = 8'h1c;
    mem[11'h0a6] = 8'h34;
    mem[11'h0a7] = 8'h1c;
    mem[11'h0a8] = 8'h9b;
    mem[11'h0a9] = 8'h1c;
    mem[11'h0aa] = 8'h33;
    mem[11'h0ab] = 8'h1b;
    mem[11'h0ac] = 8'h9d;
    mem[11'h0ad] = 8'h1c;
    mem[11'h0ae] = 8'h31;
    mem[11'h0af] = 8'h1b;
    mem[11'h0b0] = 8'h9f;
    mem[11'h0b1] = 8'h1b;
    mem[11'h0b2] = 8'h30;
    mem[11'h0b3] = 8'h86;
    mem[11'h0b4] = 8'h36;
    mem[11'h0b5] = 8'h1b;
    mem[11'h0b6] = 8'h2e;
    mem[11'h0b7] = 8'h87;
    mem[11'h0b8] = 8'h37;
    mem[11'h0b9] = 8'h1b;
    mem[11'h0ba] = 8'h2d;
    mem[11'h0bb] = 8'h87;
    mem[11'h0bc] = 8'h38;
    mem[11'h0bd] = 8'h1a;
    mem[11'h0be] = 8'h2c;
    mem[11'h0bf] = 8'h88;
    mem[11'h0c0] = 8'h39;
    mem[11'h0c1] = 8'h1a;
    mem[11'h0c2] = 8'h2a;
    mem[11'h0c3] = 8'h89;
    mem[11'h0c4] = 8'h3a;
    mem[11'h0c5] = 8'h1a;
    mem[11'h0c6] = 8'h29;
    mem[11'h0c7] = 8'h89;
    mem[11'h0c8] = 8'h3b;
    mem[11'h0c9] = 8'h19;
    mem[11'h0ca] = 8'h28;
    mem[11'h0cb] = 8'h8a;
    mem[11'h0cc] = 8'h3b;
    mem[11'h0cd] = 8'h1a;
    mem[11'h0ce] = 8'h26;
    mem[11'h0cf] = 8'h8b;
    mem[11'h0d0] = 8'h3c;
    mem[11'h0d1] = 8'h1a;
    mem[11'h0d2] = 8'h25;
    mem[11'h0d3] = 8'h8b;
    mem[11'h0d4] = 8'h3d;
    mem[11'h0d5] = 8'h19;
    mem[11'h0d6] = 8'h24;
    mem[11'h0d7] = 8'h8c;
    mem[11'h0d8] = 8'h3e;
    mem[11'h0d9] = 8'h19;
    mem[11'h0da] = 8'h23;
    mem[11'h0db] = 8'h8c;
    mem[11'h0dc] = 8'h3f;
    mem[11'h0dd] = 8'h19;
    mem[11'h0de] = 8'h21;
    mem[11'h0df] = 8'h8d;
    mem[11'h0e0] = 8'h3f;
    mem[11'h0e1] = 8'h19;
    mem[11'h0e2] = 8'h20;
    mem[11'h0e3] = 8'h8e;
    mem[11'h0e4] = 8'h40;
    mem[11'h0e5] = 8'h19;
    mem[11'h0e6] = 8'h1f;
    mem[11'h0e7] = 8'h8e;
    mem[11'h0e8] = 8'h41;
    mem[11'h0e9] = 8'h18;
    mem[11'h0ea] = 8'h1e;
    mem[11'h0eb] = 8'h8f;
    mem[11'h0ec] = 8'h41;
    mem[11'h0ed] = 8'h19;
    mem[11'h0ee] = 8'h1d;
    mem[11'h0ef] = 8'h8f;
    mem[11'h0f0] = 8'h42;
    mem[11'h0f1] = 8'h18;
    mem[11'h0f2] = 8'h1c;
    mem[11'h0f3] = 8'h90;
    mem[11'h0f4] = 8'h43;
    mem[11'h0f5] = 8'h18;
    mem[11'h0f6] = 8'h1b;
    mem[11'h0f7] = 8'h90;
    mem[11'h0f8] = 8'h43;
    mem[11'h0f9] = 8'h18;
    mem[11'h0fa] = 8'h1a;
    mem[11'h0fb] = 8'h91;
    mem[11'h0fc] = 8'h44;
    mem[11'h0fd] = 8'h18;
    mem[11'h0fe] = 8'h19;
    mem[11'h0ff] = 8'h91;
    mem[11'h100] = 8'h45;
    mem[11'h101] = 8'h17;
    mem[11'h102] = 8'h18;
    mem[11'h103] = 8'h92;
    mem[11'h104] = 8'h45;
    mem[11'h105] = 8'h18;
    mem[11'h106] = 8'h17;
    mem[11'h107] = 8'h92;
    mem[11'h108] = 8'h46;
    mem[11'h109] = 8'h17;
    mem[11'h10a] = 8'h16;
    mem[11'h10b] = 8'h93;
    mem[11'h10c] = 8'h47;
    mem[11'h10d] = 8'h17;
    mem[11'h10e] = 8'h15;
    mem[11'h10f] = 8'h93;
    mem[11'h110] = 8'h47;
    mem[11'h111] = 8'h17;
    mem[11'h112] = 8'h15;
    mem[11'h113] = 8'h93;
    mem[11'h114] = 8'h48;
    mem[11'h115] = 8'h17;
    mem[11'h116] = 8'h13;
    mem[11'h117] = 8'h94;
    mem[11'h118] = 8'h48;
    mem[11'h119] = 8'h17;
    mem[11'h11a] = 8'h13;
    mem[11'h11b] = 8'h94;
    mem[11'h11c] = 8'h49;
    mem[11'h11d] = 8'h17;
    mem[11'h11e] = 8'h11;
    mem[11'h11f] = 8'h95;
    mem[11'h120] = 8'h49;
    mem[11'h121] = 8'h17;
    mem[11'h122] = 8'h11;
    mem[11'h123] = 8'h95;
    mem[11'h124] = 8'h4a;
    mem[11'h125] = 8'h16;
    mem[11'h126] = 8'h10;
    mem[11'h127] = 8'h96;
    mem[11'h128] = 8'h4a;
    mem[11'h129] = 8'h17;
    mem[11'h12a] = 8'h0f;
    mem[11'h12b] = 8'h96;
    mem[11'h12c] = 8'h4b;
    mem[11'h12d] = 8'h16;
    mem[11'h12e] = 8'h0f;
    mem[11'h12f] = 8'h96;
    mem[11'h130] = 8'h4b;
    mem[11'h131] = 8'h16;
    mem[11'h132] = 8'h0e;
    mem[11'h133] = 8'h97;
    mem[11'h134] = 8'h4c;
    mem[11'h135] = 8'h16;
    mem[11'h136] = 8'h0d;
    mem[11'h137] = 8'h97;
    mem[11'h138] = 8'h4c;
    mem[11'h139] = 8'h16;
    mem[11'h13a] = 8'h0d;
    mem[11'h13b] = 8'h97;
    mem[11'h13c] = 8'h4d;
    mem[11'h13d] = 8'h16;
    mem[11'h13e] = 8'h0b;
    mem[11'h13f] = 8'h98;
    mem[11'h140] = 8'h4d;
    mem[11'h141] = 8'h16;
    mem[11'h142] = 8'h0b;
    mem[11'h143] = 8'h98;
    mem[11'h144] = 8'h4d;
    mem[11'h145] = 8'h16;
    mem[11'h146] = 8'h55;
    mem[11'h147] = 8'h27;
    mem[11'h148] = 8'h75;
    mem[11'h149] = 8'h16;
    mem[11'h14a] = 8'h54;
    mem[11'h14b] = 8'h27;
    mem[11'h14c] = 8'h75;
    mem[11'h14d] = 8'h16;
    mem[11'h14e] = 8'h54;
    mem[11'h14f] = 8'h27;
    mem[11'h150] = 8'h75;
    mem[11'h151] = 8'h16;
    mem[11'h152] = 8'h54;
    mem[11'h153] = 8'h27;
    mem[11'h154] = 8'h76;
    mem[11'h155] = 8'h15;
    mem[11'h156] = 8'h54;
    mem[11'h157] = 8'h27;
    mem[11'h158] = 8'h76;
    mem[11'h159] = 8'h16;
    mem[11'h15a] = 8'h53;
    mem[11'h15b] = 8'h27;
    mem[11'h15c] = 8'h77;
    mem[11'h15d] = 8'h15;
    mem[11'h15e] = 8'h53;
    mem[11'h15f] = 8'h27;
    mem[11'h160] = 8'h77;
    mem[11'h161] = 8'h15;
    mem[11'h162] = 8'h53;
    mem[11'h163] = 8'h27;
    mem[11'h164] = 8'h77;
    mem[11'h165] = 8'h16;
    mem[11'h166] = 8'h52;
    mem[11'h167] = 8'h27;
    mem[11'h168] = 8'h77;
    mem[11'h169] = 8'h16;
    mem[11'h16a] = 8'h52;
    mem[11'h16b] = 8'h27;
    mem[11'h16c] = 8'h78;
    mem[11'h16d] = 8'h15;
    mem[11'h16e] = 8'h52;
    mem[11'h16f] = 8'h27;
    mem[11'h170] = 8'h78;
    mem[11'h171] = 8'h15;
    mem[11'h172] = 8'h05;
    mem[11'h173] = 8'h15;
    mem[11'h174] = 8'h36;
    mem[11'h175] = 8'h27;
    mem[11'h176] = 8'h78;
    mem[11'h177] = 8'h15;
    mem[11'h178] = 8'h04;
    mem[11'h179] = 8'h15;
    mem[11'h17a] = 8'h37;
    mem[11'h17b] = 8'h27;
    mem[11'h17c] = 8'h79;
    mem[11'h17d] = 8'h15;
    mem[11'h17e] = 8'h03;
    mem[11'h17f] = 8'h15;
    mem[11'h180] = 8'h37;
    mem[11'h181] = 8'h27;
    mem[11'h182] = 8'h79;
    mem[11'h183] = 8'h15;
    mem[11'h184] = 8'h03;
    mem[11'h185] = 8'h15;
    mem[11'h186] = 8'h37;
    mem[11'h187] = 8'h27;
    mem[11'h188] = 8'h79;
    mem[11'h189] = 8'h15;
    mem[11'h18a] = 8'h03;
    mem[11'h18b] = 8'h15;
    mem[11'h18c] = 8'h37;
    mem[11'h18d] = 8'h27;
    mem[11'h18e] = 8'h79;
    mem[11'h18f] = 8'h15;
    mem[11'h190] = 8'h03;
    mem[11'h191] = 8'h14;
    mem[11'h192] = 8'h38;
    mem[11'h193] = 8'h27;
    mem[11'h194] = 8'h7a;
    mem[11'h195] = 8'h14;
    mem[11'h196] = 8'h02;
    mem[11'h197] = 8'h15;
    mem[11'h198] = 8'h38;
    mem[11'h199] = 8'h27;
    mem[11'h19a] = 8'h7a;
    mem[11'h19b] = 8'h15;
    mem[11'h19c] = 8'h01;
    mem[11'h19d] = 8'h15;
    mem[11'h19e] = 8'h38;
    mem[11'h19f] = 8'h27;
    mem[11'h1a0] = 8'h7a;
    mem[11'h1a1] = 8'h15;
    mem[11'h1a2] = 8'h01;
    mem[11'h1a3] = 8'h15;
    mem[11'h1a4] = 8'h38;
    mem[11'h1a5] = 8'h27;
    mem[11'h1a6] = 8'h7a;
    mem[11'h1a7] = 8'h15;
    mem[11'h1a8] = 8'h01;
    mem[11'h1a9] = 8'h15;
    mem[11'h1aa] = 8'h38;
    mem[11'h1ab] = 8'h27;
    mem[11'h1ac] = 8'h7a;
    mem[11'h1ad] = 8'h15;
    mem[11'h1ae] = 8'h01;
    mem[11'h1af] = 8'h14;
    mem[11'h1b0] = 8'h39;
    mem[11'h1b1] = 8'h27;
    mem[11'h1b2] = 8'h7b;
    mem[11'h1b3] = 8'h14;
    mem[11'h1b4] = 8'h01;
    mem[11'h1b5] = 8'h14;
    mem[11'h1b6] = 8'h39;
    mem[11'h1b7] = 8'h27;
    mem[11'h1b8] = 8'h7b;
    mem[11'h1b9] = 8'h14;
    mem[11'h1ba] = 8'h00;
    mem[11'h1bb] = 8'h15;
    mem[11'h1bc] = 8'h39;
    mem[11'h1bd] = 8'h27;
    mem[11'h1be] = 8'h7b;
    mem[11'h1bf] = 8'h2b;
    mem[11'h1c0] = 8'h39;
    mem[11'h1c1] = 8'h27;
    mem[11'h1c2] = 8'h7b;
    mem[11'h1c3] = 8'h2b;
    mem[11'h1c4] = 8'h39;
    mem[11'h1c5] = 8'h27;
    mem[11'h1c6] = 8'h7b;
    mem[11'h1c7] = 8'h2b;
    mem[11'h1c8] = 8'h39;
    mem[11'h1c9] = 8'h27;
    mem[11'h1ca] = 8'h7b;
    mem[11'h1cb] = 8'h2b;
    mem[11'h1cc] = 8'h39;
    mem[11'h1cd] = 8'h27;
    mem[11'h1ce] = 8'h7c;
    mem[11'h1cf] = 8'h29;
    mem[11'h1d0] = 8'h3a;
    mem[11'h1d1] = 8'h27;
    mem[11'h1d2] = 8'h7c;
    mem[11'h1d3] = 8'h29;
    mem[11'h1d4] = 8'h3a;
    mem[11'h1d5] = 8'h8c;
    mem[11'h1d6] = 8'h17;
    mem[11'h1d7] = 8'h29;
    mem[11'h1d8] = 8'h3a;
    mem[11'h1d9] = 8'h8c;
    mem[11'h1da] = 8'h17;
    mem[11'h1db] = 8'h29;
    mem[11'h1dc] = 8'h3a;
    mem[11'h1dd] = 8'h8c;
    mem[11'h1de] = 8'h17;
    mem[11'h1df] = 8'h29;
    mem[11'h1e0] = 8'h3a;
    mem[11'h1e1] = 8'h8c;
    mem[11'h1e2] = 8'h17;
    mem[11'h1e3] = 8'h29;
    mem[11'h1e4] = 8'h3a;
    mem[11'h1e5] = 8'h8c;
    mem[11'h1e6] = 8'h17;
    mem[11'h1e7] = 8'h29;
    mem[11'h1e8] = 8'h3a;
    mem[11'h1e9] = 8'h8c;
    mem[11'h1ea] = 8'h17;
    mem[11'h1eb] = 8'h29;
    mem[11'h1ec] = 8'h3a;
    mem[11'h1ed] = 8'h8c;
    mem[11'h1ee] = 8'h17;
    mem[11'h1ef] = 8'h29;
    mem[11'h1f0] = 8'h3a;
    mem[11'h1f1] = 8'h8c;
    mem[11'h1f2] = 8'h17;
    mem[11'h1f3] = 8'h29;
    mem[11'h1f4] = 8'h3a;
    mem[11'h1f5] = 8'h8c;
    mem[11'h1f6] = 8'h17;
    mem[11'h1f7] = 8'h29;
    mem[11'h1f8] = 8'h3a;
    mem[11'h1f9] = 8'h8c;
    mem[11'h1fa] = 8'h17;
    mem[11'h1fb] = 8'h29;
    mem[11'h1fc] = 8'h3a;
    mem[11'h1fd] = 8'h8c;
    mem[11'h1fe] = 8'h17;
    mem[11'h1ff] = 8'h29;
    mem[11'h200] = 8'h3a;
    mem[11'h201] = 8'h8c;
    mem[11'h202] = 8'h17;
    mem[11'h203] = 8'h29;
    mem[11'h204] = 8'h3a;
    mem[11'h205] = 8'h8c;
    mem[11'h206] = 8'h17;
    mem[11'h207] = 8'h29;
    mem[11'h208] = 8'h3a;
    mem[11'h209] = 8'h8c;
    mem[11'h20a] = 8'h17;
    mem[11'h20b] = 8'h29;
    mem[11'h20c] = 8'h3a;
    mem[11'h20d] = 8'h8c;
    mem[11'h20e] = 8'h17;
    mem[11'h20f] = 8'h29;
    mem[11'h210] = 8'h3a;
    mem[11'h211] = 8'h8c;
    mem[11'h212] = 8'h17;
    mem[11'h213] = 8'h29;
    mem[11'h214] = 8'h3a;
    mem[11'h215] = 8'h8c;
    mem[11'h216] = 8'h17;
    mem[11'h217] = 8'h29;
    mem[11'h218] = 8'h3a;
    mem[11'h219] = 8'h8c;
    mem[11'h21a] = 8'h17;
    mem[11'h21b] = 8'h29;
    mem[11'h21c] = 8'h3a;
    mem[11'h21d] = 8'h8c;
    mem[11'h21e] = 8'h17;
    mem[11'h21f] = 8'h29;
    mem[11'h220] = 8'h3a;
    mem[11'h221] = 8'h8c;
    mem[11'h222] = 8'h17;
    mem[11'h223] = 8'h29;
    mem[11'h224] = 8'h3a;
    mem[11'h225] = 8'h8c;
    mem[11'h226] = 8'h17;
    mem[11'h227] = 8'h29;
    mem[11'h228] = 8'h3a;
    mem[11'h229] = 8'h8c;
    mem[11'h22a] = 8'h17;
    mem[11'h22b] = 8'h29;
    mem[11'h22c] = 8'h3a;
    mem[11'h22d] = 8'h8c;
    mem[11'h22e] = 8'h17;
    mem[11'h22f] = 8'h29;
    mem[11'h230] = 8'h3a;
    mem[11'h231] = 8'h8c;
    mem[11'h232] = 8'h17;
    mem[11'h233] = 8'h29;
    mem[11'h234] = 8'h3a;
    mem[11'h235] = 8'h8c;
    mem[11'h236] = 8'h17;
    mem[11'h237] = 8'h2a;
    mem[11'h238] = 8'h39;
    mem[11'h239] = 8'h8c;
    mem[11'h23a] = 8'h17;
    mem[11'h23b] = 8'h2a;
    mem[11'h23c] = 8'h39;
    mem[11'h23d] = 8'h8c;
    mem[11'h23e] = 8'h16;
    mem[11'h23f] = 8'h2b;
    mem[11'h240] = 8'h39;
    mem[11'h241] = 8'h8c;
    mem[11'h242] = 8'h16;
    mem[11'h243] = 8'h2b;
    mem[11'h244] = 8'h39;
    mem[11'h245] = 8'h8c;
    mem[11'h246] = 8'h16;
    mem[11'h247] = 8'h15;
    mem[11'h248] = 8'h00;
    mem[11'h249] = 8'h14;
    mem[11'h24a] = 8'h39;
    mem[11'h24b] = 8'h8c;
    mem[11'h24c] = 8'h16;
    mem[11'h24d] = 8'h15;
    mem[11'h24e] = 8'h00;
    mem[11'h24f] = 8'h14;
    mem[11'h250] = 8'h39;
    mem[11'h251] = 8'h8c;
    mem[11'h252] = 8'h16;
    mem[11'h253] = 8'h14;
    mem[11'h254] = 8'h01;
    mem[11'h255] = 8'h14;
    mem[11'h256] = 8'h39;
    mem[11'h257] = 8'h8c;
    mem[11'h258] = 8'h16;
    mem[11'h259] = 8'h14;
    mem[11'h25a] = 8'h01;
    mem[11'h25b] = 8'h15;
    mem[11'h25c] = 8'h38;
    mem[11'h25d] = 8'h8c;
    mem[11'h25e] = 8'h15;
    mem[11'h25f] = 8'h15;
    mem[11'h260] = 8'h01;
    mem[11'h261] = 8'h15;
    mem[11'h262] = 8'h38;
    mem[11'h263] = 8'h8c;
    mem[11'h264] = 8'h15;
    mem[11'h265] = 8'h15;
    mem[11'h266] = 8'h01;
    mem[11'h267] = 8'h15;
    mem[11'h268] = 8'h38;
    mem[11'h269] = 8'h8c;
    mem[11'h26a] = 8'h15;
    mem[11'h26b] = 8'h15;
    mem[11'h26c] = 8'h01;
    mem[11'h26d] = 8'h15;
    mem[11'h26e] = 8'h38;
    mem[11'h26f] = 8'h8c;
    mem[11'h270] = 8'h15;
    mem[11'h271] = 8'h15;
    mem[11'h272] = 8'h02;
    mem[11'h273] = 8'h14;
    mem[11'h274] = 8'h38;
    mem[11'h275] = 8'h8c;
    mem[11'h276] = 8'h15;
    mem[11'h277] = 8'h15;
    mem[11'h278] = 8'h02;
    mem[11'h279] = 8'h15;
    mem[11'h27a] = 8'h37;
    mem[11'h27b] = 8'h27;
    mem[11'h27c] = 8'h15;
    mem[11'h27d] = 8'h27;
    mem[11'h27e] = 8'h3b;
    mem[11'h27f] = 8'h15;
    mem[11'h280] = 8'h03;
    mem[11'h281] = 8'h15;
    mem[11'h282] = 8'h37;
    mem[11'h283] = 8'h27;
    mem[11'h284] = 8'h15;
    mem[11'h285] = 8'h27;
    mem[11'h286] = 8'h3b;
    mem[11'h287] = 8'h15;
    mem[11'h288] = 8'h03;
    mem[11'h289] = 8'h15;
    mem[11'h28a] = 8'h37;
    mem[11'h28b] = 8'h27;
    mem[11'h28c] = 8'h15;
    mem[11'h28d] = 8'h27;
    mem[11'h28e] = 8'h3b;
    mem[11'h28f] = 8'h15;
    mem[11'h290] = 8'h03;
    mem[11'h291] = 8'h15;
    mem[11'h292] = 8'h37;
    mem[11'h293] = 8'h27;
    mem[11'h294] = 8'h15;
    mem[11'h295] = 8'h27;
    mem[11'h296] = 8'h3b;
    mem[11'h297] = 8'h15;
    mem[11'h298] = 8'h04;
    mem[11'h299] = 8'h15;
    mem[11'h29a] = 8'h36;
    mem[11'h29b] = 8'h27;
    mem[11'h29c] = 8'h15;
    mem[11'h29d] = 8'h27;
    mem[11'h29e] = 8'h3a;
    mem[11'h29f] = 8'h16;
    mem[11'h2a0] = 8'h04;
    mem[11'h2a1] = 8'h15;
    mem[11'h2a2] = 8'h36;
    mem[11'h2a3] = 8'h27;
    mem[11'h2a4] = 8'h15;
    mem[11'h2a5] = 8'h27;
    mem[11'h2a6] = 8'h3a;
    mem[11'h2a7] = 8'h15;
    mem[11'h2a8] = 8'h05;
    mem[11'h2a9] = 8'h15;
    mem[11'h2aa] = 8'h36;
    mem[11'h2ab] = 8'h27;
    mem[11'h2ac] = 8'h15;
    mem[11'h2ad] = 8'h27;
    mem[11'h2ae] = 8'h3a;
    mem[11'h2af] = 8'h15;
    mem[11'h2b0] = 8'h05;
    mem[11'h2b1] = 8'h16;
    mem[11'h2b2] = 8'h35;
    mem[11'h2b3] = 8'h27;
    mem[11'h2b4] = 8'h15;
    mem[11'h2b5] = 8'h27;
    mem[11'h2b6] = 8'h39;
    mem[11'h2b7] = 8'h16;
    mem[11'h2b8] = 8'h06;
    mem[11'h2b9] = 8'h15;
    mem[11'h2ba] = 8'h35;
    mem[11'h2bb] = 8'h27;
    mem[11'h2bc] = 8'h15;
    mem[11'h2bd] = 8'h27;
    mem[11'h2be] = 8'h39;
    mem[11'h2bf] = 8'h16;
    mem[11'h2c0] = 8'h06;
    mem[11'h2c1] = 8'h15;
    mem[11'h2c2] = 8'h35;
    mem[11'h2c3] = 8'h27;
    mem[11'h2c4] = 8'h15;
    mem[11'h2c5] = 8'h27;
    mem[11'h2c6] = 8'h39;
    mem[11'h2c7] = 8'h15;
    mem[11'h2c8] = 8'h07;
    mem[11'h2c9] = 8'h16;
    mem[11'h2ca] = 8'h34;
    mem[11'h2cb] = 8'h27;
    mem[11'h2cc] = 8'h15;
    mem[11'h2cd] = 8'h27;
    mem[11'h2ce] = 8'h39;
    mem[11'h2cf] = 8'h15;
    mem[11'h2d0] = 8'h07;
    mem[11'h2d1] = 8'h16;
    mem[11'h2d2] = 8'h34;
    mem[11'h2d3] = 8'h27;
    mem[11'h2d4] = 8'h15;
    mem[11'h2d5] = 8'h27;
    mem[11'h2d6] = 8'h38;
    mem[11'h2d7] = 8'h16;
    mem[11'h2d8] = 8'h08;
    mem[11'h2d9] = 8'h15;
    mem[11'h2da] = 8'h34;
    mem[11'h2db] = 8'h27;
    mem[11'h2dc] = 8'h15;
    mem[11'h2dd] = 8'h27;
    mem[11'h2de] = 8'h38;
    mem[11'h2df] = 8'h15;
    mem[11'h2e0] = 8'h09;
    mem[11'h2e1] = 8'h16;
    mem[11'h2e2] = 8'h33;
    mem[11'h2e3] = 8'h27;
    mem[11'h2e4] = 8'h15;
    mem[11'h2e5] = 8'h27;
    mem[11'h2e6] = 8'h37;
    mem[11'h2e7] = 8'h16;
    mem[11'h2e8] = 8'h09;
    mem[11'h2e9] = 8'h16;
    mem[11'h2ea] = 8'h33;
    mem[11'h2eb] = 8'h27;
    mem[11'h2ec] = 8'h15;
    mem[11'h2ed] = 8'h27;
    mem[11'h2ee] = 8'h37;
    mem[11'h2ef] = 8'h16;
    mem[11'h2f0] = 8'h0a;
    mem[11'h2f1] = 8'h15;
    mem[11'h2f2] = 8'h33;
    mem[11'h2f3] = 8'h27;
    mem[11'h2f4] = 8'h15;
    mem[11'h2f5] = 8'h27;
    mem[11'h2f6] = 8'h37;
    mem[11'h2f7] = 8'h16;
    mem[11'h2f8] = 8'h0a;
    mem[11'h2f9] = 8'h16;
    mem[11'h2fa] = 8'h32;
    mem[11'h2fb] = 8'h27;
    mem[11'h2fc] = 8'h15;
    mem[11'h2fd] = 8'h27;
    mem[11'h2fe] = 8'h36;
    mem[11'h2ff] = 8'h16;
    mem[11'h300] = 8'h0b;
    mem[11'h301] = 8'h16;
    mem[11'h302] = 8'h32;
    mem[11'h303] = 8'h27;
    mem[11'h304] = 8'h15;
    mem[11'h305] = 8'h27;
    mem[11'h306] = 8'h36;
    mem[11'h307] = 8'h16;
    mem[11'h308] = 8'h0c;
    mem[11'h309] = 8'h16;
    mem[11'h30a] = 8'h31;
    mem[11'h30b] = 8'h27;
    mem[11'h30c] = 8'h15;
    mem[11'h30d] = 8'h27;
    mem[11'h30e] = 8'h35;
    mem[11'h30f] = 8'h17;
    mem[11'h310] = 8'h0c;
    mem[11'h311] = 8'h16;
    mem[11'h312] = 8'h31;
    mem[11'h313] = 8'h27;
    mem[11'h314] = 8'h15;
    mem[11'h315] = 8'h27;
    mem[11'h316] = 8'h35;
    mem[11'h317] = 8'h16;
    mem[11'h318] = 8'h0d;
    mem[11'h319] = 8'h16;
    mem[11'h31a] = 8'h31;
    mem[11'h31b] = 8'h27;
    mem[11'h31c] = 8'h15;
    mem[11'h31d] = 8'h27;
    mem[11'h31e] = 8'h35;
    mem[11'h31f] = 8'h16;
    mem[11'h320] = 8'h0e;
    mem[11'h321] = 8'h16;
    mem[11'h322] = 8'h30;
    mem[11'h323] = 8'h27;
    mem[11'h324] = 8'h15;
    mem[11'h325] = 8'h27;
    mem[11'h326] = 8'h34;
    mem[11'h327] = 8'h17;
    mem[11'h328] = 8'h0e;
    mem[11'h329] = 8'h16;
    mem[11'h32a] = 8'h30;
    mem[11'h32b] = 8'h27;
    mem[11'h32c] = 8'h15;
    mem[11'h32d] = 8'h27;
    mem[11'h32e] = 8'h34;
    mem[11'h32f] = 8'h16;
    mem[11'h330] = 8'h0f;
    mem[11'h331] = 8'h17;
    mem[11'h332] = 8'h2f;
    mem[11'h333] = 8'h27;
    mem[11'h334] = 8'h15;
    mem[11'h335] = 8'h27;
    mem[11'h336] = 8'h33;
    mem[11'h337] = 8'h17;
    mem[11'h338] = 8'h10;
    mem[11'h339] = 8'h16;
    mem[11'h33a] = 8'h6d;
    mem[11'h33b] = 8'h27;
    mem[11'h33c] = 8'h33;
    mem[11'h33d] = 8'h16;
    mem[11'h33e] = 8'h11;
    mem[11'h33f] = 8'h17;
    mem[11'h340] = 8'h6c;
    mem[11'h341] = 8'h27;
    mem[11'h342] = 8'h32;
    mem[11'h343] = 8'h17;
    mem[11'h344] = 8'h12;
    mem[11'h345] = 8'h16;
    mem[11'h346] = 8'h6c;
    mem[11'h347] = 8'h27;
    mem[11'h348] = 8'h32;
    mem[11'h349] = 8'h17;
    mem[11'h34a] = 8'h12;
    mem[11'h34b] = 8'h17;
    mem[11'h34c] = 8'h6b;
    mem[11'h34d] = 8'h27;
    mem[11'h34e] = 8'h31;
    mem[11'h34f] = 8'h17;
    mem[11'h350] = 8'h13;
    mem[11'h351] = 8'h17;
    mem[11'h352] = 8'h6b;
    mem[11'h353] = 8'h27;
    mem[11'h354] = 8'h31;
    mem[11'h355] = 8'h17;
    mem[11'h356] = 8'h14;
    mem[11'h357] = 8'h17;
    mem[11'h358] = 8'h6a;
    mem[11'h359] = 8'h27;
    mem[11'h35a] = 8'h30;
    mem[11'h35b] = 8'h17;
    mem[11'h35c] = 8'h15;
    mem[11'h35d] = 8'h18;
    mem[11'h35e] = 8'h69;
    mem[11'h35f] = 8'h27;
    mem[11'h360] = 8'h2f;
    mem[11'h361] = 8'h18;
    mem[11'h362] = 8'h16;
    mem[11'h363] = 8'h17;
    mem[11'h364] = 8'h69;
    mem[11'h365] = 8'h27;
    mem[11'h366] = 8'h2f;
    mem[11'h367] = 8'h17;
    mem[11'h368] = 8'h17;
    mem[11'h369] = 8'h18;
    mem[11'h36a] = 8'h68;
    mem[11'h36b] = 8'h27;
    mem[11'h36c] = 8'h2e;
    mem[11'h36d] = 8'h18;
    mem[11'h36e] = 8'h18;
    mem[11'h36f] = 8'h17;
    mem[11'h370] = 8'h68;
    mem[11'h371] = 8'h27;
    mem[11'h372] = 8'h2e;
    mem[11'h373] = 8'h17;
    mem[11'h374] = 8'h19;
    mem[11'h375] = 8'h18;
    mem[11'h376] = 8'h67;
    mem[11'h377] = 8'h27;
    mem[11'h378] = 8'h2d;
    mem[11'h379] = 8'h18;
    mem[11'h37a] = 8'h1a;
    mem[11'h37b] = 8'h18;
    mem[11'h37c] = 8'h66;
    mem[11'h37d] = 8'h27;
    mem[11'h37e] = 8'h2c;
    mem[11'h37f] = 8'h18;
    mem[11'h380] = 8'h1b;
    mem[11'h381] = 8'h18;
    mem[11'h382] = 8'h66;
    mem[11'h383] = 8'h27;
    mem[11'h384] = 8'h2c;
    mem[11'h385] = 8'h18;
    mem[11'h386] = 8'h1c;
    mem[11'h387] = 8'h18;
    mem[11'h388] = 8'h65;
    mem[11'h389] = 8'h27;
    mem[11'h38a] = 8'h2b;
    mem[11'h38b] = 8'h18;
    mem[11'h38c] = 8'h1d;
    mem[11'h38d] = 8'h19;
    mem[11'h38e] = 8'h64;
    mem[11'h38f] = 8'h27;
    mem[11'h390] = 8'h2a;
    mem[11'h391] = 8'h19;
    mem[11'h392] = 8'h1e;
    mem[11'h393] = 8'h18;
    mem[11'h394] = 8'h64;
    mem[11'h395] = 8'h27;
    mem[11'h396] = 8'h2a;
    mem[11'h397] = 8'h18;
    mem[11'h398] = 8'h1f;
    mem[11'h399] = 8'h19;
    mem[11'h39a] = 8'h63;
    mem[11'h39b] = 8'h27;
    mem[11'h39c] = 8'h29;
    mem[11'h39d] = 8'h19;
    mem[11'h39e] = 8'h20;
    mem[11'h39f] = 8'h19;
    mem[11'h3a0] = 8'h62;
    mem[11'h3a1] = 8'h27;
    mem[11'h3a2] = 8'h28;
    mem[11'h3a3] = 8'h19;
    mem[11'h3a4] = 8'h22;
    mem[11'h3a5] = 8'h19;
    mem[11'h3a6] = 8'h61;
    mem[11'h3a7] = 8'h27;
    mem[11'h3a8] = 8'h28;
    mem[11'h3a9] = 8'h19;
    mem[11'h3aa] = 8'h22;
    mem[11'h3ab] = 8'h19;
    mem[11'h3ac] = 8'h61;
    mem[11'h3ad] = 8'h27;
    mem[11'h3ae] = 8'h27;
    mem[11'h3af] = 8'h19;
    mem[11'h3b0] = 8'h24;
    mem[11'h3b1] = 8'h19;
    mem[11'h3b2] = 8'h60;
    mem[11'h3b3] = 8'h27;
    mem[11'h3b4] = 8'h26;
    mem[11'h3b5] = 8'h19;
    mem[11'h3b6] = 8'h25;
    mem[11'h3b7] = 8'h1a;
    mem[11'h3b8] = 8'h5f;
    mem[11'h3b9] = 8'h27;
    mem[11'h3ba] = 8'h25;
    mem[11'h3bb] = 8'h1a;
    mem[11'h3bc] = 8'h26;
    mem[11'h3bd] = 8'h1a;
    mem[11'h3be] = 8'h5e;
    mem[11'h3bf] = 8'h27;
    mem[11'h3c0] = 8'h24;
    mem[11'h3c1] = 8'h1a;
    mem[11'h3c2] = 8'h28;
    mem[11'h3c3] = 8'h1a;
    mem[11'h3c4] = 8'h5d;
    mem[11'h3c5] = 8'h27;
    mem[11'h3c6] = 8'h24;
    mem[11'h3c7] = 8'h19;
    mem[11'h3c8] = 8'h29;
    mem[11'h3c9] = 8'h1a;
    mem[11'h3ca] = 8'h5d;
    mem[11'h3cb] = 8'h27;
    mem[11'h3cc] = 8'h23;
    mem[11'h3cd] = 8'h1a;
    mem[11'h3ce] = 8'h2a;
    mem[11'h3cf] = 8'h1a;
    mem[11'h3d0] = 8'h5c;
    mem[11'h3d1] = 8'h27;
    mem[11'h3d2] = 8'h22;
    mem[11'h3d3] = 8'h1a;
    mem[11'h3d4] = 8'h2c;
    mem[11'h3d5] = 8'h1a;
    mem[11'h3d6] = 8'h5b;
    mem[11'h3d7] = 8'h27;
    mem[11'h3d8] = 8'h21;
    mem[11'h3d9] = 8'h1a;
    mem[11'h3da] = 8'h2d;
    mem[11'h3db] = 8'h1b;
    mem[11'h3dc] = 8'h5a;
    mem[11'h3dd] = 8'h27;
    mem[11'h3de] = 8'h20;
    mem[11'h3df] = 8'h1b;
    mem[11'h3e0] = 8'h2e;
    mem[11'h3e1] = 8'h1b;
    mem[11'h3e2] = 8'h59;
    mem[11'h3e3] = 8'h27;
    mem[11'h3e4] = 8'h1f;
    mem[11'h3e5] = 8'h1b;
    mem[11'h3e6] = 8'h30;
    mem[11'h3e7] = 8'h1b;
    mem[11'h3e8] = 8'h58;
    mem[11'h3e9] = 8'h27;
    mem[11'h3ea] = 8'h1e;
    mem[11'h3eb] = 8'h1b;
    mem[11'h3ec] = 8'h32;
    mem[11'h3ed] = 8'h1b;
    mem[11'h3ee] = 8'h57;
    mem[11'h3ef] = 8'h27;
    mem[11'h3f0] = 8'h1d;
    mem[11'h3f1] = 8'h1c;
    mem[11'h3f2] = 8'h32;
    mem[11'h3f3] = 8'h1c;
    mem[11'h3f4] = 8'h56;
    mem[11'h3f5] = 8'h27;
    mem[11'h3f6] = 8'h1c;
    mem[11'h3f7] = 8'h1c;
    mem[11'h3f8] = 8'h34;
    mem[11'h3f9] = 8'h1c;
    mem[11'h3fa] = 8'h55;
    mem[11'h3fb] = 8'h27;
    mem[11'h3fc] = 8'h1b;
    mem[11'h3fd] = 8'h1c;
    mem[11'h3fe] = 8'h36;
    mem[11'h3ff] = 8'h1c;
    mem[11'h400] = 8'h54;
    mem[11'h401] = 8'h27;
    mem[11'h402] = 8'h1a;
    mem[11'h403] = 8'h1c;
    mem[11'h404] = 8'h38;
    mem[11'h405] = 8'h1c;
    mem[11'h406] = 8'h53;
    mem[11'h407] = 8'h27;
    mem[11'h408] = 8'h19;
    mem[11'h409] = 8'h1d;
    mem[11'h40a] = 8'h38;
    mem[11'h40b] = 8'h1d;
    mem[11'h40c] = 8'h52;
    mem[11'h40d] = 8'h27;
    mem[11'h40e] = 8'h18;
    mem[11'h40f] = 8'h1d;
    mem[11'h410] = 8'h3a;
    mem[11'h411] = 8'h1e;
    mem[11'h412] = 8'h50;
    mem[11'h413] = 8'h27;
    mem[11'h414] = 8'h16;
    mem[11'h415] = 8'h1e;
    mem[11'h416] = 8'h3c;
    mem[11'h417] = 8'h1e;
    mem[11'h418] = 8'h4f;
    mem[11'h419] = 8'h27;
    mem[11'h41a] = 8'h15;
    mem[11'h41b] = 8'h1e;
    mem[11'h41c] = 8'h3e;
    mem[11'h41d] = 8'h1e;
    mem[11'h41e] = 8'h4e;
    mem[11'h41f] = 8'h27;
    mem[11'h420] = 8'h14;
    mem[11'h421] = 8'h1e;
    mem[11'h422] = 8'h40;
    mem[11'h423] = 8'h1e;
    mem[11'h424] = 8'h4d;
    mem[11'h425] = 8'h27;
    mem[11'h426] = 8'h13;
    mem[11'h427] = 8'h1e;
    mem[11'h428] = 8'h42;
    mem[11'h429] = 8'h1f;
    mem[11'h42a] = 8'h4b;
    mem[11'h42b] = 8'h27;
    mem[11'h42c] = 8'h11;
    mem[11'h42d] = 8'h1f;
    mem[11'h42e] = 8'h44;
    mem[11'h42f] = 8'h1f;
    mem[11'h430] = 8'h4a;
    mem[11'h431] = 8'h27;
    mem[11'h432] = 8'h10;
    mem[11'h433] = 8'h20;
    mem[11'h434] = 8'h45;
    mem[11'h435] = 8'h1f;
    mem[11'h436] = 8'h49;
    mem[11'h437] = 8'h27;
    mem[11'h438] = 8'h0f;
    mem[11'h439] = 8'h20;
    mem[11'h43a] = 8'h47;
    mem[11'h43b] = 8'h20;
    mem[11'h43c] = 8'h47;
    mem[11'h43d] = 8'h27;
    mem[11'h43e] = 8'h0d;
    mem[11'h43f] = 8'h21;
    mem[11'h440] = 8'h49;
    mem[11'h441] = 8'h20;
    mem[11'h442] = 8'h46;
    mem[11'h443] = 8'h27;
    mem[11'h444] = 8'h0c;
    mem[11'h445] = 8'h21;
    mem[11'h446] = 8'h4a;
    mem[11'h447] = 8'h22;
    mem[11'h448] = 8'h44;
    mem[11'h449] = 8'h27;
    mem[11'h44a] = 8'h0a;
    mem[11'h44b] = 8'h22;
    mem[11'h44c] = 8'h4d;
    mem[11'h44d] = 8'h21;
    mem[11'h44e] = 8'h43;
    mem[11'h44f] = 8'h27;
    mem[11'h450] = 8'h0a;
    mem[11'h451] = 8'h21;
    mem[11'h452] = 8'h4f;
    mem[11'h453] = 8'h22;
    mem[11'h454] = 8'h41;
    mem[11'h455] = 8'h27;
    mem[11'h456] = 8'h0a;
    mem[11'h457] = 8'h20;
    mem[11'h458] = 8'h51;
    mem[11'h459] = 8'h23;
    mem[11'h45a] = 8'h3f;
    mem[11'h45b] = 8'h27;
    mem[11'h45c] = 8'h0a;
    mem[11'h45d] = 8'h1f;
    mem[11'h45e] = 8'h53;
    mem[11'h45f] = 8'h23;
    mem[11'h460] = 8'h3e;
    mem[11'h461] = 8'h27;
    mem[11'h462] = 8'h0a;
    mem[11'h463] = 8'h1e;
    mem[11'h464] = 8'h55;
    mem[11'h465] = 8'h24;
    mem[11'h466] = 8'h3c;
    mem[11'h467] = 8'h27;
    mem[11'h468] = 8'h0a;
    mem[11'h469] = 8'h1c;
    mem[11'h46a] = 8'h58;
    mem[11'h46b] = 8'h25;
    mem[11'h46c] = 8'h3a;
    mem[11'h46d] = 8'h27;
    mem[11'h46e] = 8'h0a;
    mem[11'h46f] = 8'h1b;
    mem[11'h470] = 8'h5a;
    mem[11'h471] = 8'h26;
    mem[11'h472] = 8'h38;
    mem[11'h473] = 8'h27;
    mem[11'h474] = 8'h0a;
    mem[11'h475] = 8'h1a;
    mem[11'h476] = 8'h5c;
    mem[11'h477] = 8'h28;
    mem[11'h478] = 8'h35;
    mem[11'h479] = 8'h27;
    mem[11'h47a] = 8'h0a;
    mem[11'h47b] = 8'h19;
    mem[11'h47c] = 8'h5e;
    mem[11'h47d] = 8'h29;
    mem[11'h47e] = 8'h33;
    mem[11'h47f] = 8'h27;
    mem[11'h480] = 8'h0a;
    mem[11'h481] = 8'h18;
    mem[11'h482] = 8'h61;
    mem[11'h483] = 8'h29;
    mem[11'h484] = 8'h31;
    mem[11'h485] = 8'h27;
    mem[11'h486] = 8'h0a;
    mem[11'h487] = 8'h17;
    mem[11'h488] = 8'h63;
    mem[11'h489] = 8'h2b;
    mem[11'h48a] = 8'h2e;
    mem[11'h48b] = 8'h27;
    mem[11'h48c] = 8'h0a;
    mem[11'h48d] = 8'h15;
    mem[11'h48e] = 8'h66;
    mem[11'h48f] = 8'h2d;
    mem[11'h490] = 8'h2b;
    mem[11'h491] = 8'h27;
    mem[11'h492] = 8'h0a;
    mem[11'h493] = 8'h14;
    mem[11'h494] = 8'h69;
    mem[11'h495] = 8'h2e;
    mem[11'h496] = 8'h28;
    mem[11'h497] = 8'h27;
    mem[11'h498] = 8'h0a;
    mem[11'h499] = 8'h13;
    mem[11'h49a] = 8'h6b;
    mem[11'h49b] = 8'h31;
    mem[11'h49c] = 8'h24;
    mem[11'h49d] = 8'h27;
    mem[11'h49e] = 8'h0a;
    mem[11'h49f] = 8'h11;
    mem[11'h4a0] = 8'h6e;
    mem[11'h4a1] = 8'h34;
    mem[11'h4a2] = 8'h20;
    mem[11'h4a3] = 8'h27;
    mem[11'h4a4] = 8'h0a;
    mem[11'h4a5] = 8'h10;
    mem[11'h4a6] = 8'h71;
    mem[11'h4a7] = 8'h37;
    mem[11'h4a8] = 8'h1b;
    mem[11'h4a9] = 8'h27;
    mem[11'h4aa] = 8'h0a;
    mem[11'h4ab] = 8'h0e;
    mem[11'h4ac] = 8'h74;
    mem[11'h4ad] = 8'h3c;
    mem[11'h4ae] = 8'h15;
    mem[11'h4af] = 8'h27;
    mem[11'h4b0] = 8'h0a;
    mem[11'h4b1] = 8'h0d;
    mem[11'h4b2] = 8'h77;
    mem[11'h4b3] = 8'h78;
    mem[11'h4b4] = 8'h0a;
    mem[11'h4b5] = 8'h0b;
    mem[11'h4b6] = 8'h7a;
    mem[11'h4b7] = 8'h77;
    mem[11'h4b8] = 8'h0a;
    mem[11'h4b9] = 8'h0a;
    mem[11'h4ba] = 8'h7d;
    mem[11'h4bb] = 8'h75;
    mem[11'h4bc] = 8'h0a;
    mem[11'h4bd] = 8'h08;
    mem[11'h4be] = 8'h81;
    mem[11'h4bf] = 8'h73;
    mem[11'h4c0] = 8'h0a;
    mem[11'h4c1] = 8'h06;
    mem[11'h4c2] = 8'h85;
    mem[11'h4c3] = 8'h71;
    mem[11'h4c4] = 8'h0a;
    mem[11'h4c5] = 8'h05;
    mem[11'h4c6] = 8'h87;
    mem[11'h4c7] = 8'h70;
    mem[11'h4c8] = 8'h0a;
    mem[11'h4c9] = 8'h03;
    mem[11'h4ca] = 8'h8b;
    mem[11'h4cb] = 8'h6e;
    mem[11'h4cc] = 8'h0a;
    mem[11'h4cd] = 8'h01;
    mem[11'h4ce] = 8'h8f;
    mem[11'h4cf] = 8'h6c;
    mem[11'h4d0] = 8'h9e;
    mem[11'h4d1] = 8'h6a;
    mem[11'h4d2] = 8'ha0;
    mem[11'h4d3] = 8'h68;
    mem[11'h4d4] = 8'ha3;
    mem[11'h4d5] = 8'h65;
    mem[11'h4d6] = 8'ha5;
    mem[11'h4d7] = 8'h63;
    mem[11'h4d8] = 8'ha7;
    mem[11'h4d9] = 8'h61;
    mem[11'h4da] = 8'haa;
    mem[11'h4db] = 8'h5b;
    mem[11'h4dc] = 8'hb0;
    mem[11'h4dd] = 8'h55;
    mem[11'h4de] = 8'hb6;
    mem[11'h4df] = 8'h4f;
    mem[11'h4e0] = 8'hbc;
    mem[11'h4e1] = 8'h49;
    mem[11'h4e2] = 8'hc3;
    mem[11'h4e3] = 8'h41;
    mem[11'h4e4] = 8'hcb;
    mem[11'h4e5] = 8'h39;
    mem[11'h4e6] = 8'hd5;
    mem[11'h4e7] = 8'h2e;
    mem[11'h4e8] = 8'he0;
    mem[11'h4e9] = 8'h21;
    mem[11'h4ea] = 8'hff;
    mem[11'h4eb] = 8'hff;
  end
  assign len = mem[addr];
endmodule

