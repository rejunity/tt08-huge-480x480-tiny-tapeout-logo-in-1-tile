/*
 * Copyright (c) 2024 Tiny Tapeout LTD
 * SPDX-License-Identifier: Apache-2.0
 * Author: Renaldas Zioma
 */

`default_nettype none

parameter LOGO_SIZE = 128;  // Size of the logo in pixels
parameter DISPLAY_WIDTH = 640;  // VGA display width
parameter DISPLAY_HEIGHT = 480;  // VGA display height

`define COLOR_WHITE 3'd7

module tt_um_rejunity_vga_logo (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // VGA signals
  wire hsync;
  wire vsync;
  reg [1:0] R;
  reg [1:0] G;
  reg [1:0] B;
  wire video_active;
  wire [9:0] pix_x;
  wire [9:0] pix_y;


  // TinyVGA PMOD
  assign uo_out  = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

  // Unused outputs assigned to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in[7:1], uio_in};

  hvsync_generator vga_sync_gen (
      .clk(clk),
      .reset(~rst_n),
      .hsync(hsync),
      .vsync(vsync),
      .display_on(video_active),
      .hpos(pix_x),
      .vpos(pix_y)
  );

  reg pixel_value;

  // bitmap_rom rom1 (
  //     .x(pix_x[6:0]),
  //     .y(pix_y[6:0]),
  //     .pixel(pixel_value)
  // );

  reg [11:0] addr;
  reg [7:0] len;
  bitmap_rom_rle rom2 (
    .addr(addr),
    .len(len)
  );

  assign {R, G, B } = video_active*pixel_value*6'b11_11_00;

  // increase couner every frame (vsync happens once per frame)
  reg [11:0] counter;
  always @(posedge clk) begin
    if (~rst_n) begin
      counter <= 0;
    end else begin
      if (vsync) begin
        addr <= 0;
        counter <= 0;
        pixel_value <= 0;
      end else if (pix_x < 272 && pix_y < 267) begin
        if (counter >= len) begin
          addr <= addr + 1;
          counter <= 0;
          pixel_value <= ~pixel_value;
        end else
          counter <= counter + 1;
      end
    end
  end  

endmodule

// --------------------------------------------------------

module bitmap_rom_rle (
    input wire [11:0] addr,
    output wire [7:0] len
);

  reg [7:0] mem[1329:0];
  initial begin
    mem[12'h000] = 8'h87;
    mem[12'h001] = 8'h01;
    mem[12'h002] = 8'hfd;
    mem[12'h003] = 8'h21;
    mem[12'h004] = 8'he7;
    mem[12'h005] = 8'h2d;
    mem[12'h006] = 8'hdc;
    mem[12'h007] = 8'h38;
    mem[12'h008] = 8'hd1;
    mem[12'h009] = 8'h41;
    mem[12'h00a] = 8'hca;
    mem[12'h00b] = 8'h48;
    mem[12'h00c] = 8'hc2;
    mem[12'h00d] = 8'h4f;
    mem[12'h00e] = 8'hbc;
    mem[12'h00f] = 8'h55;
    mem[12'h010] = 8'hb6;
    mem[12'h011] = 8'h5b;
    mem[12'h012] = 8'hb0;
    mem[12'h013] = 8'h61;
    mem[12'h014] = 8'hab;
    mem[12'h015] = 8'h65;
    mem[12'h016] = 8'ha7;
    mem[12'h017] = 8'h69;
    mem[12'h018] = 8'ha2;
    mem[12'h019] = 8'h6f;
    mem[12'h01a] = 8'h9d;
    mem[12'h01b] = 8'h73;
    mem[12'h01c] = 8'h99;
    mem[12'h01d] = 8'h77;
    mem[12'h01e] = 8'h95;
    mem[12'h01f] = 8'h7b;
    mem[12'h020] = 8'h91;
    mem[12'h021] = 8'h7f;
    mem[12'h022] = 8'h8e;
    mem[12'h023] = 8'h82;
    mem[12'h024] = 8'h8a;
    mem[12'h025] = 8'h85;
    mem[12'h026] = 8'h87;
    mem[12'h027] = 8'h89;
    mem[12'h028] = 8'h84;
    mem[12'h029] = 8'h8c;
    mem[12'h02a] = 8'h80;
    mem[12'h02b] = 8'h8f;
    mem[12'h02c] = 8'h7d;
    mem[12'h02d] = 8'h3c;
    mem[12'h02e] = 8'h19;
    mem[12'h02f] = 8'h3c;
    mem[12'h030] = 8'h7a;
    mem[12'h031] = 8'h37;
    mem[12'h032] = 8'h25;
    mem[12'h033] = 8'h37;
    mem[12'h034] = 8'h77;
    mem[12'h035] = 8'h34;
    mem[12'h036] = 8'h2f;
    mem[12'h037] = 8'h34;
    mem[12'h038] = 8'h74;
    mem[12'h039] = 8'h31;
    mem[12'h03a] = 8'h38;
    mem[12'h03b] = 8'h30;
    mem[12'h03c] = 8'h72;
    mem[12'h03d] = 8'h2e;
    mem[12'h03e] = 8'h3f;
    mem[12'h03f] = 8'h2e;
    mem[12'h040] = 8'h6f;
    mem[12'h041] = 8'h2d;
    mem[12'h042] = 8'h45;
    mem[12'h043] = 8'h2d;
    mem[12'h044] = 8'h6c;
    mem[12'h045] = 8'h2b;
    mem[12'h046] = 8'h4b;
    mem[12'h047] = 8'h2b;
    mem[12'h048] = 8'h6a;
    mem[12'h049] = 8'h29;
    mem[12'h04a] = 8'h51;
    mem[12'h04b] = 8'h29;
    mem[12'h04c] = 8'h68;
    mem[12'h04d] = 8'h28;
    mem[12'h04e] = 8'h55;
    mem[12'h04f] = 8'h29;
    mem[12'h050] = 8'h64;
    mem[12'h051] = 8'h28;
    mem[12'h052] = 8'h59;
    mem[12'h053] = 8'h28;
    mem[12'h054] = 8'h62;
    mem[12'h055] = 8'h27;
    mem[12'h056] = 8'h5e;
    mem[12'h057] = 8'h26;
    mem[12'h058] = 8'h60;
    mem[12'h059] = 8'h25;
    mem[12'h05a] = 8'h63;
    mem[12'h05b] = 8'h25;
    mem[12'h05c] = 8'h5e;
    mem[12'h05d] = 8'h24;
    mem[12'h05e] = 8'h67;
    mem[12'h05f] = 8'h24;
    mem[12'h060] = 8'h5c;
    mem[12'h061] = 8'h24;
    mem[12'h062] = 8'h6a;
    mem[12'h063] = 8'h23;
    mem[12'h064] = 8'h5a;
    mem[12'h065] = 8'h23;
    mem[12'h066] = 8'h6d;
    mem[12'h067] = 8'h23;
    mem[12'h068] = 8'h58;
    mem[12'h069] = 8'h22;
    mem[12'h06a] = 8'h71;
    mem[12'h06b] = 8'h23;
    mem[12'h06c] = 8'h55;
    mem[12'h06d] = 8'h21;
    mem[12'h06e] = 8'h75;
    mem[12'h06f] = 8'h22;
    mem[12'h070] = 8'h53;
    mem[12'h071] = 8'h21;
    mem[12'h072] = 8'h77;
    mem[12'h073] = 8'h22;
    mem[12'h074] = 8'h51;
    mem[12'h075] = 8'h20;
    mem[12'h076] = 8'h7b;
    mem[12'h077] = 8'h21;
    mem[12'h078] = 8'h4f;
    mem[12'h079] = 8'h20;
    mem[12'h07a] = 8'h7d;
    mem[12'h07b] = 8'h21;
    mem[12'h07c] = 8'h4d;
    mem[12'h07d] = 8'h1f;
    mem[12'h07e] = 8'h81;
    mem[12'h07f] = 8'h1f;
    mem[12'h080] = 8'h4c;
    mem[12'h081] = 8'h1f;
    mem[12'h082] = 8'h83;
    mem[12'h083] = 8'h1f;
    mem[12'h084] = 8'h4a;
    mem[12'h085] = 8'h1f;
    mem[12'h086] = 8'h85;
    mem[12'h087] = 8'h1f;
    mem[12'h088] = 8'h48;
    mem[12'h089] = 8'h1e;
    mem[12'h08a] = 8'h89;
    mem[12'h08b] = 8'h1e;
    mem[12'h08c] = 8'h46;
    mem[12'h08d] = 8'h1e;
    mem[12'h08e] = 8'h8b;
    mem[12'h08f] = 8'h1e;
    mem[12'h090] = 8'h44;
    mem[12'h091] = 8'h1e;
    mem[12'h092] = 8'h8d;
    mem[12'h093] = 8'h1e;
    mem[12'h094] = 8'h42;
    mem[12'h095] = 8'h1e;
    mem[12'h096] = 8'h8f;
    mem[12'h097] = 8'h1e;
    mem[12'h098] = 8'h40;
    mem[12'h099] = 8'h1d;
    mem[12'h09a] = 8'h93;
    mem[12'h09b] = 8'h1d;
    mem[12'h09c] = 8'h3f;
    mem[12'h09d] = 8'h1c;
    mem[12'h09e] = 8'h95;
    mem[12'h09f] = 8'h1c;
    mem[12'h0a0] = 8'h3e;
    mem[12'h0a1] = 8'h1c;
    mem[12'h0a2] = 8'h97;
    mem[12'h0a3] = 8'h1c;
    mem[12'h0a4] = 8'h3c;
    mem[12'h0a5] = 8'h1c;
    mem[12'h0a6] = 8'h99;
    mem[12'h0a7] = 8'h1c;
    mem[12'h0a8] = 8'h3a;
    mem[12'h0a9] = 8'h1c;
    mem[12'h0aa] = 8'h9b;
    mem[12'h0ab] = 8'h1c;
    mem[12'h0ac] = 8'h39;
    mem[12'h0ad] = 8'h1b;
    mem[12'h0ae] = 8'h9d;
    mem[12'h0af] = 8'h1c;
    mem[12'h0b0] = 8'h37;
    mem[12'h0b1] = 8'h1b;
    mem[12'h0b2] = 8'h9f;
    mem[12'h0b3] = 8'h1b;
    mem[12'h0b4] = 8'h36;
    mem[12'h0b5] = 8'h86;
    mem[12'h0b6] = 8'h36;
    mem[12'h0b7] = 8'h1b;
    mem[12'h0b8] = 8'h34;
    mem[12'h0b9] = 8'h87;
    mem[12'h0ba] = 8'h37;
    mem[12'h0bb] = 8'h1b;
    mem[12'h0bc] = 8'h33;
    mem[12'h0bd] = 8'h87;
    mem[12'h0be] = 8'h38;
    mem[12'h0bf] = 8'h1a;
    mem[12'h0c0] = 8'h32;
    mem[12'h0c1] = 8'h88;
    mem[12'h0c2] = 8'h39;
    mem[12'h0c3] = 8'h1a;
    mem[12'h0c4] = 8'h30;
    mem[12'h0c5] = 8'h89;
    mem[12'h0c6] = 8'h3a;
    mem[12'h0c7] = 8'h1a;
    mem[12'h0c8] = 8'h2f;
    mem[12'h0c9] = 8'h89;
    mem[12'h0ca] = 8'h3a;
    mem[12'h0cb] = 8'h1a;
    mem[12'h0cc] = 8'h2e;
    mem[12'h0cd] = 8'h8a;
    mem[12'h0ce] = 8'h3b;
    mem[12'h0cf] = 8'h1a;
    mem[12'h0d0] = 8'h2c;
    mem[12'h0d1] = 8'h8b;
    mem[12'h0d2] = 8'h3c;
    mem[12'h0d3] = 8'h1a;
    mem[12'h0d4] = 8'h2b;
    mem[12'h0d5] = 8'h8b;
    mem[12'h0d6] = 8'h3d;
    mem[12'h0d7] = 8'h19;
    mem[12'h0d8] = 8'h2a;
    mem[12'h0d9] = 8'h8c;
    mem[12'h0da] = 8'h3e;
    mem[12'h0db] = 8'h19;
    mem[12'h0dc] = 8'h29;
    mem[12'h0dd] = 8'h8c;
    mem[12'h0de] = 8'h3e;
    mem[12'h0df] = 8'h19;
    mem[12'h0e0] = 8'h28;
    mem[12'h0e1] = 8'h8d;
    mem[12'h0e2] = 8'h3f;
    mem[12'h0e3] = 8'h19;
    mem[12'h0e4] = 8'h27;
    mem[12'h0e5] = 8'h8d;
    mem[12'h0e6] = 8'h40;
    mem[12'h0e7] = 8'h19;
    mem[12'h0e8] = 8'h25;
    mem[12'h0e9] = 8'h8e;
    mem[12'h0ea] = 8'h41;
    mem[12'h0eb] = 8'h18;
    mem[12'h0ec] = 8'h24;
    mem[12'h0ed] = 8'h8f;
    mem[12'h0ee] = 8'h41;
    mem[12'h0ef] = 8'h19;
    mem[12'h0f0] = 8'h23;
    mem[12'h0f1] = 8'h8f;
    mem[12'h0f2] = 8'h42;
    mem[12'h0f3] = 8'h18;
    mem[12'h0f4] = 8'h22;
    mem[12'h0f5] = 8'h90;
    mem[12'h0f6] = 8'h43;
    mem[12'h0f7] = 8'h18;
    mem[12'h0f8] = 8'h21;
    mem[12'h0f9] = 8'h90;
    mem[12'h0fa] = 8'h43;
    mem[12'h0fb] = 8'h18;
    mem[12'h0fc] = 8'h20;
    mem[12'h0fd] = 8'h91;
    mem[12'h0fe] = 8'h44;
    mem[12'h0ff] = 8'h18;
    mem[12'h100] = 8'h1f;
    mem[12'h101] = 8'h91;
    mem[12'h102] = 8'h45;
    mem[12'h103] = 8'h17;
    mem[12'h104] = 8'h1e;
    mem[12'h105] = 8'h92;
    mem[12'h106] = 8'h45;
    mem[12'h107] = 8'h18;
    mem[12'h108] = 8'h1d;
    mem[12'h109] = 8'h92;
    mem[12'h10a] = 8'h46;
    mem[12'h10b] = 8'h17;
    mem[12'h10c] = 8'h1c;
    mem[12'h10d] = 8'h93;
    mem[12'h10e] = 8'h46;
    mem[12'h10f] = 8'h18;
    mem[12'h110] = 8'h1b;
    mem[12'h111] = 8'h93;
    mem[12'h112] = 8'h47;
    mem[12'h113] = 8'h17;
    mem[12'h114] = 8'h1b;
    mem[12'h115] = 8'h93;
    mem[12'h116] = 8'h48;
    mem[12'h117] = 8'h17;
    mem[12'h118] = 8'h19;
    mem[12'h119] = 8'h94;
    mem[12'h11a] = 8'h48;
    mem[12'h11b] = 8'h17;
    mem[12'h11c] = 8'h19;
    mem[12'h11d] = 8'h94;
    mem[12'h11e] = 8'h49;
    mem[12'h11f] = 8'h16;
    mem[12'h120] = 8'h18;
    mem[12'h121] = 8'h95;
    mem[12'h122] = 8'h49;
    mem[12'h123] = 8'h17;
    mem[12'h124] = 8'h17;
    mem[12'h125] = 8'h95;
    mem[12'h126] = 8'h4a;
    mem[12'h127] = 8'h16;
    mem[12'h128] = 8'h16;
    mem[12'h129] = 8'h96;
    mem[12'h12a] = 8'h4a;
    mem[12'h12b] = 8'h17;
    mem[12'h12c] = 8'h15;
    mem[12'h12d] = 8'h96;
    mem[12'h12e] = 8'h4b;
    mem[12'h12f] = 8'h16;
    mem[12'h130] = 8'h15;
    mem[12'h131] = 8'h96;
    mem[12'h132] = 8'h4b;
    mem[12'h133] = 8'h16;
    mem[12'h134] = 8'h14;
    mem[12'h135] = 8'h97;
    mem[12'h136] = 8'h4c;
    mem[12'h137] = 8'h16;
    mem[12'h138] = 8'h13;
    mem[12'h139] = 8'h97;
    mem[12'h13a] = 8'h4c;
    mem[12'h13b] = 8'h16;
    mem[12'h13c] = 8'h13;
    mem[12'h13d] = 8'h97;
    mem[12'h13e] = 8'h4c;
    mem[12'h13f] = 8'h16;
    mem[12'h140] = 8'h12;
    mem[12'h141] = 8'h98;
    mem[12'h142] = 8'h4d;
    mem[12'h143] = 8'h16;
    mem[12'h144] = 8'h11;
    mem[12'h145] = 8'h98;
    mem[12'h146] = 8'h4d;
    mem[12'h147] = 8'h16;
    mem[12'h148] = 8'h5b;
    mem[12'h149] = 8'h27;
    mem[12'h14a] = 8'h75;
    mem[12'h14b] = 8'h16;
    mem[12'h14c] = 8'h5a;
    mem[12'h14d] = 8'h27;
    mem[12'h14e] = 8'h75;
    mem[12'h14f] = 8'h16;
    mem[12'h150] = 8'h5a;
    mem[12'h151] = 8'h27;
    mem[12'h152] = 8'h75;
    mem[12'h153] = 8'h16;
    mem[12'h154] = 8'h5a;
    mem[12'h155] = 8'h27;
    mem[12'h156] = 8'h76;
    mem[12'h157] = 8'h15;
    mem[12'h158] = 8'h5a;
    mem[12'h159] = 8'h27;
    mem[12'h15a] = 8'h76;
    mem[12'h15b] = 8'h16;
    mem[12'h15c] = 8'h59;
    mem[12'h15d] = 8'h27;
    mem[12'h15e] = 8'h76;
    mem[12'h15f] = 8'h16;
    mem[12'h160] = 8'h59;
    mem[12'h161] = 8'h27;
    mem[12'h162] = 8'h77;
    mem[12'h163] = 8'h15;
    mem[12'h164] = 8'h59;
    mem[12'h165] = 8'h27;
    mem[12'h166] = 8'h77;
    mem[12'h167] = 8'h16;
    mem[12'h168] = 8'h58;
    mem[12'h169] = 8'h27;
    mem[12'h16a] = 8'h77;
    mem[12'h16b] = 8'h16;
    mem[12'h16c] = 8'h58;
    mem[12'h16d] = 8'h27;
    mem[12'h16e] = 8'h78;
    mem[12'h16f] = 8'h15;
    mem[12'h170] = 8'h58;
    mem[12'h171] = 8'h27;
    mem[12'h172] = 8'h78;
    mem[12'h173] = 8'h15;
    mem[12'h174] = 8'h0b;
    mem[12'h175] = 8'h15;
    mem[12'h176] = 8'h36;
    mem[12'h177] = 8'h27;
    mem[12'h178] = 8'h78;
    mem[12'h179] = 8'h15;
    mem[12'h17a] = 8'h0a;
    mem[12'h17b] = 8'h16;
    mem[12'h17c] = 8'h36;
    mem[12'h17d] = 8'h27;
    mem[12'h17e] = 8'h79;
    mem[12'h17f] = 8'h15;
    mem[12'h180] = 8'h09;
    mem[12'h181] = 8'h15;
    mem[12'h182] = 8'h37;
    mem[12'h183] = 8'h27;
    mem[12'h184] = 8'h79;
    mem[12'h185] = 8'h15;
    mem[12'h186] = 8'h09;
    mem[12'h187] = 8'h15;
    mem[12'h188] = 8'h37;
    mem[12'h189] = 8'h27;
    mem[12'h18a] = 8'h79;
    mem[12'h18b] = 8'h15;
    mem[12'h18c] = 8'h09;
    mem[12'h18d] = 8'h15;
    mem[12'h18e] = 8'h37;
    mem[12'h18f] = 8'h27;
    mem[12'h190] = 8'h79;
    mem[12'h191] = 8'h15;
    mem[12'h192] = 8'h09;
    mem[12'h193] = 8'h15;
    mem[12'h194] = 8'h37;
    mem[12'h195] = 8'h27;
    mem[12'h196] = 8'h7a;
    mem[12'h197] = 8'h14;
    mem[12'h198] = 8'h08;
    mem[12'h199] = 8'h15;
    mem[12'h19a] = 8'h38;
    mem[12'h19b] = 8'h27;
    mem[12'h19c] = 8'h7a;
    mem[12'h19d] = 8'h15;
    mem[12'h19e] = 8'h07;
    mem[12'h19f] = 8'h15;
    mem[12'h1a0] = 8'h38;
    mem[12'h1a1] = 8'h27;
    mem[12'h1a2] = 8'h7a;
    mem[12'h1a3] = 8'h15;
    mem[12'h1a4] = 8'h07;
    mem[12'h1a5] = 8'h15;
    mem[12'h1a6] = 8'h38;
    mem[12'h1a7] = 8'h27;
    mem[12'h1a8] = 8'h7a;
    mem[12'h1a9] = 8'h15;
    mem[12'h1aa] = 8'h07;
    mem[12'h1ab] = 8'h15;
    mem[12'h1ac] = 8'h38;
    mem[12'h1ad] = 8'h27;
    mem[12'h1ae] = 8'h7a;
    mem[12'h1af] = 8'h15;
    mem[12'h1b0] = 8'h07;
    mem[12'h1b1] = 8'h15;
    mem[12'h1b2] = 8'h38;
    mem[12'h1b3] = 8'h27;
    mem[12'h1b4] = 8'h7b;
    mem[12'h1b5] = 8'h14;
    mem[12'h1b6] = 8'h07;
    mem[12'h1b7] = 8'h14;
    mem[12'h1b8] = 8'h39;
    mem[12'h1b9] = 8'h27;
    mem[12'h1ba] = 8'h7b;
    mem[12'h1bb] = 8'h14;
    mem[12'h1bc] = 8'h06;
    mem[12'h1bd] = 8'h15;
    mem[12'h1be] = 8'h39;
    mem[12'h1bf] = 8'h27;
    mem[12'h1c0] = 8'h7b;
    mem[12'h1c1] = 8'h15;
    mem[12'h1c2] = 8'h05;
    mem[12'h1c3] = 8'h15;
    mem[12'h1c4] = 8'h39;
    mem[12'h1c5] = 8'h27;
    mem[12'h1c6] = 8'h7b;
    mem[12'h1c7] = 8'h15;
    mem[12'h1c8] = 8'h05;
    mem[12'h1c9] = 8'h15;
    mem[12'h1ca] = 8'h39;
    mem[12'h1cb] = 8'h27;
    mem[12'h1cc] = 8'h7b;
    mem[12'h1cd] = 8'h15;
    mem[12'h1ce] = 8'h05;
    mem[12'h1cf] = 8'h15;
    mem[12'h1d0] = 8'h39;
    mem[12'h1d1] = 8'h27;
    mem[12'h1d2] = 8'h7b;
    mem[12'h1d3] = 8'h15;
    mem[12'h1d4] = 8'h05;
    mem[12'h1d5] = 8'h15;
    mem[12'h1d6] = 8'h39;
    mem[12'h1d7] = 8'h27;
    mem[12'h1d8] = 8'h7b;
    mem[12'h1d9] = 8'h15;
    mem[12'h1da] = 8'h05;
    mem[12'h1db] = 8'h14;
    mem[12'h1dc] = 8'h3a;
    mem[12'h1dd] = 8'h27;
    mem[12'h1de] = 8'h7c;
    mem[12'h1df] = 8'h14;
    mem[12'h1e0] = 8'h05;
    mem[12'h1e1] = 8'h14;
    mem[12'h1e2] = 8'h3a;
    mem[12'h1e3] = 8'h8c;
    mem[12'h1e4] = 8'h17;
    mem[12'h1e5] = 8'h14;
    mem[12'h1e6] = 8'h05;
    mem[12'h1e7] = 8'h14;
    mem[12'h1e8] = 8'h3a;
    mem[12'h1e9] = 8'h8c;
    mem[12'h1ea] = 8'h17;
    mem[12'h1eb] = 8'h14;
    mem[12'h1ec] = 8'h05;
    mem[12'h1ed] = 8'h14;
    mem[12'h1ee] = 8'h3a;
    mem[12'h1ef] = 8'h8c;
    mem[12'h1f0] = 8'h17;
    mem[12'h1f1] = 8'h14;
    mem[12'h1f2] = 8'h05;
    mem[12'h1f3] = 8'h14;
    mem[12'h1f4] = 8'h3a;
    mem[12'h1f5] = 8'h8c;
    mem[12'h1f6] = 8'h17;
    mem[12'h1f7] = 8'h14;
    mem[12'h1f8] = 8'h05;
    mem[12'h1f9] = 8'h14;
    mem[12'h1fa] = 8'h3a;
    mem[12'h1fb] = 8'h8c;
    mem[12'h1fc] = 8'h17;
    mem[12'h1fd] = 8'h15;
    mem[12'h1fe] = 8'h04;
    mem[12'h1ff] = 8'h14;
    mem[12'h200] = 8'h3a;
    mem[12'h201] = 8'h8c;
    mem[12'h202] = 8'h17;
    mem[12'h203] = 8'h15;
    mem[12'h204] = 8'h04;
    mem[12'h205] = 8'h14;
    mem[12'h206] = 8'h3a;
    mem[12'h207] = 8'h8c;
    mem[12'h208] = 8'h17;
    mem[12'h209] = 8'h15;
    mem[12'h20a] = 8'h03;
    mem[12'h20b] = 8'h15;
    mem[12'h20c] = 8'h3a;
    mem[12'h20d] = 8'h8c;
    mem[12'h20e] = 8'h17;
    mem[12'h20f] = 8'h15;
    mem[12'h210] = 8'h03;
    mem[12'h211] = 8'h15;
    mem[12'h212] = 8'h3a;
    mem[12'h213] = 8'h8c;
    mem[12'h214] = 8'h17;
    mem[12'h215] = 8'h15;
    mem[12'h216] = 8'h03;
    mem[12'h217] = 8'h15;
    mem[12'h218] = 8'h3a;
    mem[12'h219] = 8'h8c;
    mem[12'h21a] = 8'h17;
    mem[12'h21b] = 8'h15;
    mem[12'h21c] = 8'h03;
    mem[12'h21d] = 8'h15;
    mem[12'h21e] = 8'h3a;
    mem[12'h21f] = 8'h8c;
    mem[12'h220] = 8'h17;
    mem[12'h221] = 8'h15;
    mem[12'h222] = 8'h03;
    mem[12'h223] = 8'h15;
    mem[12'h224] = 8'h3a;
    mem[12'h225] = 8'h8c;
    mem[12'h226] = 8'h17;
    mem[12'h227] = 8'h15;
    mem[12'h228] = 8'h03;
    mem[12'h229] = 8'h15;
    mem[12'h22a] = 8'h3a;
    mem[12'h22b] = 8'h8c;
    mem[12'h22c] = 8'h17;
    mem[12'h22d] = 8'h15;
    mem[12'h22e] = 8'h03;
    mem[12'h22f] = 8'h15;
    mem[12'h230] = 8'h3a;
    mem[12'h231] = 8'h8c;
    mem[12'h232] = 8'h17;
    mem[12'h233] = 8'h15;
    mem[12'h234] = 8'h03;
    mem[12'h235] = 8'h15;
    mem[12'h236] = 8'h3a;
    mem[12'h237] = 8'h8c;
    mem[12'h238] = 8'h17;
    mem[12'h239] = 8'h15;
    mem[12'h23a] = 8'h03;
    mem[12'h23b] = 8'h15;
    mem[12'h23c] = 8'h3a;
    mem[12'h23d] = 8'h8c;
    mem[12'h23e] = 8'h17;
    mem[12'h23f] = 8'h15;
    mem[12'h240] = 8'h03;
    mem[12'h241] = 8'h15;
    mem[12'h242] = 8'h3a;
    mem[12'h243] = 8'h8c;
    mem[12'h244] = 8'h17;
    mem[12'h245] = 8'h15;
    mem[12'h246] = 8'h03;
    mem[12'h247] = 8'h15;
    mem[12'h248] = 8'h3a;
    mem[12'h249] = 8'h8c;
    mem[12'h24a] = 8'h17;
    mem[12'h24b] = 8'h15;
    mem[12'h24c] = 8'h04;
    mem[12'h24d] = 8'h14;
    mem[12'h24e] = 8'h3a;
    mem[12'h24f] = 8'h8c;
    mem[12'h250] = 8'h17;
    mem[12'h251] = 8'h15;
    mem[12'h252] = 8'h04;
    mem[12'h253] = 8'h14;
    mem[12'h254] = 8'h3a;
    mem[12'h255] = 8'h8c;
    mem[12'h256] = 8'h17;
    mem[12'h257] = 8'h15;
    mem[12'h258] = 8'h04;
    mem[12'h259] = 8'h14;
    mem[12'h25a] = 8'h3a;
    mem[12'h25b] = 8'h8c;
    mem[12'h25c] = 8'h17;
    mem[12'h25d] = 8'h14;
    mem[12'h25e] = 8'h05;
    mem[12'h25f] = 8'h14;
    mem[12'h260] = 8'h3a;
    mem[12'h261] = 8'h8c;
    mem[12'h262] = 8'h17;
    mem[12'h263] = 8'h14;
    mem[12'h264] = 8'h05;
    mem[12'h265] = 8'h14;
    mem[12'h266] = 8'h3a;
    mem[12'h267] = 8'h8c;
    mem[12'h268] = 8'h17;
    mem[12'h269] = 8'h14;
    mem[12'h26a] = 8'h05;
    mem[12'h26b] = 8'h14;
    mem[12'h26c] = 8'h3a;
    mem[12'h26d] = 8'h8c;
    mem[12'h26e] = 8'h17;
    mem[12'h26f] = 8'h14;
    mem[12'h270] = 8'h05;
    mem[12'h271] = 8'h14;
    mem[12'h272] = 8'h3a;
    mem[12'h273] = 8'h8c;
    mem[12'h274] = 8'h17;
    mem[12'h275] = 8'h14;
    mem[12'h276] = 8'h05;
    mem[12'h277] = 8'h15;
    mem[12'h278] = 8'h39;
    mem[12'h279] = 8'h8c;
    mem[12'h27a] = 8'h17;
    mem[12'h27b] = 8'h14;
    mem[12'h27c] = 8'h05;
    mem[12'h27d] = 8'h15;
    mem[12'h27e] = 8'h39;
    mem[12'h27f] = 8'h8c;
    mem[12'h280] = 8'h16;
    mem[12'h281] = 8'h15;
    mem[12'h282] = 8'h05;
    mem[12'h283] = 8'h15;
    mem[12'h284] = 8'h39;
    mem[12'h285] = 8'h8c;
    mem[12'h286] = 8'h16;
    mem[12'h287] = 8'h15;
    mem[12'h288] = 8'h05;
    mem[12'h289] = 8'h15;
    mem[12'h28a] = 8'h39;
    mem[12'h28b] = 8'h8c;
    mem[12'h28c] = 8'h16;
    mem[12'h28d] = 8'h15;
    mem[12'h28e] = 8'h05;
    mem[12'h28f] = 8'h15;
    mem[12'h290] = 8'h39;
    mem[12'h291] = 8'h8c;
    mem[12'h292] = 8'h16;
    mem[12'h293] = 8'h15;
    mem[12'h294] = 8'h06;
    mem[12'h295] = 8'h14;
    mem[12'h296] = 8'h39;
    mem[12'h297] = 8'h8c;
    mem[12'h298] = 8'h16;
    mem[12'h299] = 8'h15;
    mem[12'h29a] = 8'h06;
    mem[12'h29b] = 8'h14;
    mem[12'h29c] = 8'h39;
    mem[12'h29d] = 8'h8c;
    mem[12'h29e] = 8'h16;
    mem[12'h29f] = 8'h14;
    mem[12'h2a0] = 8'h07;
    mem[12'h2a1] = 8'h15;
    mem[12'h2a2] = 8'h38;
    mem[12'h2a3] = 8'h8c;
    mem[12'h2a4] = 8'h15;
    mem[12'h2a5] = 8'h15;
    mem[12'h2a6] = 8'h07;
    mem[12'h2a7] = 8'h15;
    mem[12'h2a8] = 8'h38;
    mem[12'h2a9] = 8'h8c;
    mem[12'h2aa] = 8'h15;
    mem[12'h2ab] = 8'h15;
    mem[12'h2ac] = 8'h07;
    mem[12'h2ad] = 8'h15;
    mem[12'h2ae] = 8'h38;
    mem[12'h2af] = 8'h8c;
    mem[12'h2b0] = 8'h15;
    mem[12'h2b1] = 8'h15;
    mem[12'h2b2] = 8'h07;
    mem[12'h2b3] = 8'h15;
    mem[12'h2b4] = 8'h38;
    mem[12'h2b5] = 8'h8c;
    mem[12'h2b6] = 8'h15;
    mem[12'h2b7] = 8'h15;
    mem[12'h2b8] = 8'h08;
    mem[12'h2b9] = 8'h14;
    mem[12'h2ba] = 8'h38;
    mem[12'h2bb] = 8'h8c;
    mem[12'h2bc] = 8'h15;
    mem[12'h2bd] = 8'h15;
    mem[12'h2be] = 8'h08;
    mem[12'h2bf] = 8'h15;
    mem[12'h2c0] = 8'h37;
    mem[12'h2c1] = 8'h27;
    mem[12'h2c2] = 8'h15;
    mem[12'h2c3] = 8'h27;
    mem[12'h2c4] = 8'h3b;
    mem[12'h2c5] = 8'h15;
    mem[12'h2c6] = 8'h09;
    mem[12'h2c7] = 8'h15;
    mem[12'h2c8] = 8'h37;
    mem[12'h2c9] = 8'h27;
    mem[12'h2ca] = 8'h15;
    mem[12'h2cb] = 8'h27;
    mem[12'h2cc] = 8'h3b;
    mem[12'h2cd] = 8'h15;
    mem[12'h2ce] = 8'h09;
    mem[12'h2cf] = 8'h15;
    mem[12'h2d0] = 8'h37;
    mem[12'h2d1] = 8'h27;
    mem[12'h2d2] = 8'h15;
    mem[12'h2d3] = 8'h27;
    mem[12'h2d4] = 8'h3b;
    mem[12'h2d5] = 8'h15;
    mem[12'h2d6] = 8'h09;
    mem[12'h2d7] = 8'h15;
    mem[12'h2d8] = 8'h37;
    mem[12'h2d9] = 8'h27;
    mem[12'h2da] = 8'h15;
    mem[12'h2db] = 8'h27;
    mem[12'h2dc] = 8'h3b;
    mem[12'h2dd] = 8'h15;
    mem[12'h2de] = 8'h0a;
    mem[12'h2df] = 8'h15;
    mem[12'h2e0] = 8'h36;
    mem[12'h2e1] = 8'h27;
    mem[12'h2e2] = 8'h15;
    mem[12'h2e3] = 8'h27;
    mem[12'h2e4] = 8'h3a;
    mem[12'h2e5] = 8'h16;
    mem[12'h2e6] = 8'h0a;
    mem[12'h2e7] = 8'h15;
    mem[12'h2e8] = 8'h36;
    mem[12'h2e9] = 8'h27;
    mem[12'h2ea] = 8'h15;
    mem[12'h2eb] = 8'h27;
    mem[12'h2ec] = 8'h3a;
    mem[12'h2ed] = 8'h15;
    mem[12'h2ee] = 8'h0b;
    mem[12'h2ef] = 8'h15;
    mem[12'h2f0] = 8'h36;
    mem[12'h2f1] = 8'h27;
    mem[12'h2f2] = 8'h15;
    mem[12'h2f3] = 8'h27;
    mem[12'h2f4] = 8'h3a;
    mem[12'h2f5] = 8'h15;
    mem[12'h2f6] = 8'h0b;
    mem[12'h2f7] = 8'h16;
    mem[12'h2f8] = 8'h35;
    mem[12'h2f9] = 8'h27;
    mem[12'h2fa] = 8'h15;
    mem[12'h2fb] = 8'h27;
    mem[12'h2fc] = 8'h39;
    mem[12'h2fd] = 8'h16;
    mem[12'h2fe] = 8'h0c;
    mem[12'h2ff] = 8'h15;
    mem[12'h300] = 8'h35;
    mem[12'h301] = 8'h27;
    mem[12'h302] = 8'h15;
    mem[12'h303] = 8'h27;
    mem[12'h304] = 8'h39;
    mem[12'h305] = 8'h16;
    mem[12'h306] = 8'h0c;
    mem[12'h307] = 8'h15;
    mem[12'h308] = 8'h35;
    mem[12'h309] = 8'h27;
    mem[12'h30a] = 8'h15;
    mem[12'h30b] = 8'h27;
    mem[12'h30c] = 8'h39;
    mem[12'h30d] = 8'h15;
    mem[12'h30e] = 8'h0d;
    mem[12'h30f] = 8'h16;
    mem[12'h310] = 8'h34;
    mem[12'h311] = 8'h27;
    mem[12'h312] = 8'h15;
    mem[12'h313] = 8'h27;
    mem[12'h314] = 8'h39;
    mem[12'h315] = 8'h15;
    mem[12'h316] = 8'h0d;
    mem[12'h317] = 8'h16;
    mem[12'h318] = 8'h34;
    mem[12'h319] = 8'h27;
    mem[12'h31a] = 8'h15;
    mem[12'h31b] = 8'h27;
    mem[12'h31c] = 8'h38;
    mem[12'h31d] = 8'h16;
    mem[12'h31e] = 8'h0e;
    mem[12'h31f] = 8'h15;
    mem[12'h320] = 8'h34;
    mem[12'h321] = 8'h27;
    mem[12'h322] = 8'h15;
    mem[12'h323] = 8'h27;
    mem[12'h324] = 8'h38;
    mem[12'h325] = 8'h16;
    mem[12'h326] = 8'h0e;
    mem[12'h327] = 8'h16;
    mem[12'h328] = 8'h33;
    mem[12'h329] = 8'h27;
    mem[12'h32a] = 8'h15;
    mem[12'h32b] = 8'h27;
    mem[12'h32c] = 8'h37;
    mem[12'h32d] = 8'h16;
    mem[12'h32e] = 8'h0f;
    mem[12'h32f] = 8'h16;
    mem[12'h330] = 8'h33;
    mem[12'h331] = 8'h27;
    mem[12'h332] = 8'h15;
    mem[12'h333] = 8'h27;
    mem[12'h334] = 8'h37;
    mem[12'h335] = 8'h16;
    mem[12'h336] = 8'h10;
    mem[12'h337] = 8'h15;
    mem[12'h338] = 8'h33;
    mem[12'h339] = 8'h27;
    mem[12'h33a] = 8'h15;
    mem[12'h33b] = 8'h27;
    mem[12'h33c] = 8'h37;
    mem[12'h33d] = 8'h16;
    mem[12'h33e] = 8'h10;
    mem[12'h33f] = 8'h16;
    mem[12'h340] = 8'h32;
    mem[12'h341] = 8'h27;
    mem[12'h342] = 8'h15;
    mem[12'h343] = 8'h27;
    mem[12'h344] = 8'h36;
    mem[12'h345] = 8'h16;
    mem[12'h346] = 8'h11;
    mem[12'h347] = 8'h16;
    mem[12'h348] = 8'h32;
    mem[12'h349] = 8'h27;
    mem[12'h34a] = 8'h15;
    mem[12'h34b] = 8'h27;
    mem[12'h34c] = 8'h36;
    mem[12'h34d] = 8'h16;
    mem[12'h34e] = 8'h12;
    mem[12'h34f] = 8'h16;
    mem[12'h350] = 8'h31;
    mem[12'h351] = 8'h27;
    mem[12'h352] = 8'h15;
    mem[12'h353] = 8'h27;
    mem[12'h354] = 8'h35;
    mem[12'h355] = 8'h17;
    mem[12'h356] = 8'h12;
    mem[12'h357] = 8'h16;
    mem[12'h358] = 8'h31;
    mem[12'h359] = 8'h27;
    mem[12'h35a] = 8'h15;
    mem[12'h35b] = 8'h27;
    mem[12'h35c] = 8'h35;
    mem[12'h35d] = 8'h16;
    mem[12'h35e] = 8'h13;
    mem[12'h35f] = 8'h16;
    mem[12'h360] = 8'h31;
    mem[12'h361] = 8'h27;
    mem[12'h362] = 8'h15;
    mem[12'h363] = 8'h27;
    mem[12'h364] = 8'h35;
    mem[12'h365] = 8'h16;
    mem[12'h366] = 8'h14;
    mem[12'h367] = 8'h16;
    mem[12'h368] = 8'h30;
    mem[12'h369] = 8'h27;
    mem[12'h36a] = 8'h15;
    mem[12'h36b] = 8'h27;
    mem[12'h36c] = 8'h34;
    mem[12'h36d] = 8'h17;
    mem[12'h36e] = 8'h14;
    mem[12'h36f] = 8'h16;
    mem[12'h370] = 8'h30;
    mem[12'h371] = 8'h27;
    mem[12'h372] = 8'h15;
    mem[12'h373] = 8'h27;
    mem[12'h374] = 8'h34;
    mem[12'h375] = 8'h16;
    mem[12'h376] = 8'h15;
    mem[12'h377] = 8'h17;
    mem[12'h378] = 8'h2f;
    mem[12'h379] = 8'h27;
    mem[12'h37a] = 8'h15;
    mem[12'h37b] = 8'h27;
    mem[12'h37c] = 8'h33;
    mem[12'h37d] = 8'h17;
    mem[12'h37e] = 8'h16;
    mem[12'h37f] = 8'h16;
    mem[12'h380] = 8'h6d;
    mem[12'h381] = 8'h27;
    mem[12'h382] = 8'h33;
    mem[12'h383] = 8'h16;
    mem[12'h384] = 8'h17;
    mem[12'h385] = 8'h17;
    mem[12'h386] = 8'h6c;
    mem[12'h387] = 8'h27;
    mem[12'h388] = 8'h32;
    mem[12'h389] = 8'h17;
    mem[12'h38a] = 8'h18;
    mem[12'h38b] = 8'h16;
    mem[12'h38c] = 8'h6c;
    mem[12'h38d] = 8'h27;
    mem[12'h38e] = 8'h32;
    mem[12'h38f] = 8'h17;
    mem[12'h390] = 8'h18;
    mem[12'h391] = 8'h17;
    mem[12'h392] = 8'h6b;
    mem[12'h393] = 8'h27;
    mem[12'h394] = 8'h31;
    mem[12'h395] = 8'h17;
    mem[12'h396] = 8'h19;
    mem[12'h397] = 8'h17;
    mem[12'h398] = 8'h6b;
    mem[12'h399] = 8'h27;
    mem[12'h39a] = 8'h31;
    mem[12'h39b] = 8'h17;
    mem[12'h39c] = 8'h1a;
    mem[12'h39d] = 8'h17;
    mem[12'h39e] = 8'h6a;
    mem[12'h39f] = 8'h27;
    mem[12'h3a0] = 8'h30;
    mem[12'h3a1] = 8'h17;
    mem[12'h3a2] = 8'h1b;
    mem[12'h3a3] = 8'h18;
    mem[12'h3a4] = 8'h69;
    mem[12'h3a5] = 8'h27;
    mem[12'h3a6] = 8'h30;
    mem[12'h3a7] = 8'h17;
    mem[12'h3a8] = 8'h1c;
    mem[12'h3a9] = 8'h17;
    mem[12'h3aa] = 8'h69;
    mem[12'h3ab] = 8'h27;
    mem[12'h3ac] = 8'h2f;
    mem[12'h3ad] = 8'h17;
    mem[12'h3ae] = 8'h1d;
    mem[12'h3af] = 8'h18;
    mem[12'h3b0] = 8'h68;
    mem[12'h3b1] = 8'h27;
    mem[12'h3b2] = 8'h2e;
    mem[12'h3b3] = 8'h18;
    mem[12'h3b4] = 8'h1e;
    mem[12'h3b5] = 8'h17;
    mem[12'h3b6] = 8'h68;
    mem[12'h3b7] = 8'h27;
    mem[12'h3b8] = 8'h2e;
    mem[12'h3b9] = 8'h17;
    mem[12'h3ba] = 8'h1f;
    mem[12'h3bb] = 8'h18;
    mem[12'h3bc] = 8'h67;
    mem[12'h3bd] = 8'h27;
    mem[12'h3be] = 8'h2d;
    mem[12'h3bf] = 8'h18;
    mem[12'h3c0] = 8'h20;
    mem[12'h3c1] = 8'h18;
    mem[12'h3c2] = 8'h66;
    mem[12'h3c3] = 8'h27;
    mem[12'h3c4] = 8'h2d;
    mem[12'h3c5] = 8'h17;
    mem[12'h3c6] = 8'h21;
    mem[12'h3c7] = 8'h18;
    mem[12'h3c8] = 8'h66;
    mem[12'h3c9] = 8'h27;
    mem[12'h3ca] = 8'h2c;
    mem[12'h3cb] = 8'h18;
    mem[12'h3cc] = 8'h22;
    mem[12'h3cd] = 8'h18;
    mem[12'h3ce] = 8'h65;
    mem[12'h3cf] = 8'h27;
    mem[12'h3d0] = 8'h2b;
    mem[12'h3d1] = 8'h18;
    mem[12'h3d2] = 8'h23;
    mem[12'h3d3] = 8'h19;
    mem[12'h3d4] = 8'h64;
    mem[12'h3d5] = 8'h27;
    mem[12'h3d6] = 8'h2a;
    mem[12'h3d7] = 8'h19;
    mem[12'h3d8] = 8'h24;
    mem[12'h3d9] = 8'h18;
    mem[12'h3da] = 8'h64;
    mem[12'h3db] = 8'h27;
    mem[12'h3dc] = 8'h2a;
    mem[12'h3dd] = 8'h18;
    mem[12'h3de] = 8'h25;
    mem[12'h3df] = 8'h19;
    mem[12'h3e0] = 8'h63;
    mem[12'h3e1] = 8'h27;
    mem[12'h3e2] = 8'h29;
    mem[12'h3e3] = 8'h19;
    mem[12'h3e4] = 8'h26;
    mem[12'h3e5] = 8'h19;
    mem[12'h3e6] = 8'h62;
    mem[12'h3e7] = 8'h27;
    mem[12'h3e8] = 8'h28;
    mem[12'h3e9] = 8'h19;
    mem[12'h3ea] = 8'h28;
    mem[12'h3eb] = 8'h18;
    mem[12'h3ec] = 8'h62;
    mem[12'h3ed] = 8'h27;
    mem[12'h3ee] = 8'h28;
    mem[12'h3ef] = 8'h19;
    mem[12'h3f0] = 8'h28;
    mem[12'h3f1] = 8'h19;
    mem[12'h3f2] = 8'h61;
    mem[12'h3f3] = 8'h27;
    mem[12'h3f4] = 8'h27;
    mem[12'h3f5] = 8'h19;
    mem[12'h3f6] = 8'h2a;
    mem[12'h3f7] = 8'h19;
    mem[12'h3f8] = 8'h60;
    mem[12'h3f9] = 8'h27;
    mem[12'h3fa] = 8'h26;
    mem[12'h3fb] = 8'h19;
    mem[12'h3fc] = 8'h2b;
    mem[12'h3fd] = 8'h1a;
    mem[12'h3fe] = 8'h5f;
    mem[12'h3ff] = 8'h27;
    mem[12'h400] = 8'h25;
    mem[12'h401] = 8'h1a;
    mem[12'h402] = 8'h2c;
    mem[12'h403] = 8'h1a;
    mem[12'h404] = 8'h5e;
    mem[12'h405] = 8'h27;
    mem[12'h406] = 8'h24;
    mem[12'h407] = 8'h1a;
    mem[12'h408] = 8'h2e;
    mem[12'h409] = 8'h19;
    mem[12'h40a] = 8'h5e;
    mem[12'h40b] = 8'h27;
    mem[12'h40c] = 8'h24;
    mem[12'h40d] = 8'h1a;
    mem[12'h40e] = 8'h2e;
    mem[12'h40f] = 8'h1a;
    mem[12'h410] = 8'h5d;
    mem[12'h411] = 8'h27;
    mem[12'h412] = 8'h23;
    mem[12'h413] = 8'h1a;
    mem[12'h414] = 8'h30;
    mem[12'h415] = 8'h1a;
    mem[12'h416] = 8'h5c;
    mem[12'h417] = 8'h27;
    mem[12'h418] = 8'h22;
    mem[12'h419] = 8'h1a;
    mem[12'h41a] = 8'h32;
    mem[12'h41b] = 8'h1a;
    mem[12'h41c] = 8'h5b;
    mem[12'h41d] = 8'h27;
    mem[12'h41e] = 8'h21;
    mem[12'h41f] = 8'h1b;
    mem[12'h420] = 8'h32;
    mem[12'h421] = 8'h1b;
    mem[12'h422] = 8'h5a;
    mem[12'h423] = 8'h27;
    mem[12'h424] = 8'h20;
    mem[12'h425] = 8'h1b;
    mem[12'h426] = 8'h34;
    mem[12'h427] = 8'h1b;
    mem[12'h428] = 8'h59;
    mem[12'h429] = 8'h27;
    mem[12'h42a] = 8'h1f;
    mem[12'h42b] = 8'h1b;
    mem[12'h42c] = 8'h36;
    mem[12'h42d] = 8'h1b;
    mem[12'h42e] = 8'h58;
    mem[12'h42f] = 8'h27;
    mem[12'h430] = 8'h1e;
    mem[12'h431] = 8'h1b;
    mem[12'h432] = 8'h37;
    mem[12'h433] = 8'h1c;
    mem[12'h434] = 8'h57;
    mem[12'h435] = 8'h27;
    mem[12'h436] = 8'h1d;
    mem[12'h437] = 8'h1c;
    mem[12'h438] = 8'h38;
    mem[12'h439] = 8'h1c;
    mem[12'h43a] = 8'h56;
    mem[12'h43b] = 8'h27;
    mem[12'h43c] = 8'h1c;
    mem[12'h43d] = 8'h1c;
    mem[12'h43e] = 8'h3a;
    mem[12'h43f] = 8'h1c;
    mem[12'h440] = 8'h55;
    mem[12'h441] = 8'h27;
    mem[12'h442] = 8'h1b;
    mem[12'h443] = 8'h1c;
    mem[12'h444] = 8'h3c;
    mem[12'h445] = 8'h1c;
    mem[12'h446] = 8'h54;
    mem[12'h447] = 8'h27;
    mem[12'h448] = 8'h1a;
    mem[12'h449] = 8'h1c;
    mem[12'h44a] = 8'h3e;
    mem[12'h44b] = 8'h1c;
    mem[12'h44c] = 8'h53;
    mem[12'h44d] = 8'h27;
    mem[12'h44e] = 8'h19;
    mem[12'h44f] = 8'h1d;
    mem[12'h450] = 8'h3e;
    mem[12'h451] = 8'h1d;
    mem[12'h452] = 8'h52;
    mem[12'h453] = 8'h27;
    mem[12'h454] = 8'h18;
    mem[12'h455] = 8'h1d;
    mem[12'h456] = 8'h40;
    mem[12'h457] = 8'h1d;
    mem[12'h458] = 8'h51;
    mem[12'h459] = 8'h27;
    mem[12'h45a] = 8'h17;
    mem[12'h45b] = 8'h1d;
    mem[12'h45c] = 8'h42;
    mem[12'h45d] = 8'h1e;
    mem[12'h45e] = 8'h4f;
    mem[12'h45f] = 8'h27;
    mem[12'h460] = 8'h15;
    mem[12'h461] = 8'h1e;
    mem[12'h462] = 8'h44;
    mem[12'h463] = 8'h1e;
    mem[12'h464] = 8'h4e;
    mem[12'h465] = 8'h27;
    mem[12'h466] = 8'h14;
    mem[12'h467] = 8'h1e;
    mem[12'h468] = 8'h46;
    mem[12'h469] = 8'h1e;
    mem[12'h46a] = 8'h4d;
    mem[12'h46b] = 8'h27;
    mem[12'h46c] = 8'h13;
    mem[12'h46d] = 8'h1e;
    mem[12'h46e] = 8'h48;
    mem[12'h46f] = 8'h1e;
    mem[12'h470] = 8'h4c;
    mem[12'h471] = 8'h27;
    mem[12'h472] = 8'h12;
    mem[12'h473] = 8'h1e;
    mem[12'h474] = 8'h49;
    mem[12'h475] = 8'h20;
    mem[12'h476] = 8'h4a;
    mem[12'h477] = 8'h27;
    mem[12'h478] = 8'h10;
    mem[12'h479] = 8'h20;
    mem[12'h47a] = 8'h4a;
    mem[12'h47b] = 8'h20;
    mem[12'h47c] = 8'h49;
    mem[12'h47d] = 8'h27;
    mem[12'h47e] = 8'h0f;
    mem[12'h47f] = 8'h20;
    mem[12'h480] = 8'h4c;
    mem[12'h481] = 8'h21;
    mem[12'h482] = 8'h47;
    mem[12'h483] = 8'h27;
    mem[12'h484] = 8'h0d;
    mem[12'h485] = 8'h21;
    mem[12'h486] = 8'h4e;
    mem[12'h487] = 8'h21;
    mem[12'h488] = 8'h46;
    mem[12'h489] = 8'h27;
    mem[12'h48a] = 8'h0c;
    mem[12'h48b] = 8'h21;
    mem[12'h48c] = 8'h50;
    mem[12'h48d] = 8'h22;
    mem[12'h48e] = 8'h44;
    mem[12'h48f] = 8'h27;
    mem[12'h490] = 8'h0b;
    mem[12'h491] = 8'h21;
    mem[12'h492] = 8'h52;
    mem[12'h493] = 8'h22;
    mem[12'h494] = 8'h43;
    mem[12'h495] = 8'h27;
    mem[12'h496] = 8'h0a;
    mem[12'h497] = 8'h21;
    mem[12'h498] = 8'h54;
    mem[12'h499] = 8'h23;
    mem[12'h49a] = 8'h41;
    mem[12'h49b] = 8'h27;
    mem[12'h49c] = 8'h0a;
    mem[12'h49d] = 8'h20;
    mem[12'h49e] = 8'h56;
    mem[12'h49f] = 8'h24;
    mem[12'h4a0] = 8'h3f;
    mem[12'h4a1] = 8'h27;
    mem[12'h4a2] = 8'h0a;
    mem[12'h4a3] = 8'h1f;
    mem[12'h4a4] = 8'h58;
    mem[12'h4a5] = 8'h24;
    mem[12'h4a6] = 8'h3e;
    mem[12'h4a7] = 8'h27;
    mem[12'h4a8] = 8'h0a;
    mem[12'h4a9] = 8'h1e;
    mem[12'h4aa] = 8'h5b;
    mem[12'h4ab] = 8'h24;
    mem[12'h4ac] = 8'h3c;
    mem[12'h4ad] = 8'h27;
    mem[12'h4ae] = 8'h0a;
    mem[12'h4af] = 8'h1d;
    mem[12'h4b0] = 8'h5d;
    mem[12'h4b1] = 8'h25;
    mem[12'h4b2] = 8'h3a;
    mem[12'h4b3] = 8'h27;
    mem[12'h4b4] = 8'h0a;
    mem[12'h4b5] = 8'h1b;
    mem[12'h4b6] = 8'h60;
    mem[12'h4b7] = 8'h26;
    mem[12'h4b8] = 8'h38;
    mem[12'h4b9] = 8'h27;
    mem[12'h4ba] = 8'h0a;
    mem[12'h4bb] = 8'h1a;
    mem[12'h4bc] = 8'h62;
    mem[12'h4bd] = 8'h27;
    mem[12'h4be] = 8'h36;
    mem[12'h4bf] = 8'h27;
    mem[12'h4c0] = 8'h0a;
    mem[12'h4c1] = 8'h19;
    mem[12'h4c2] = 8'h64;
    mem[12'h4c3] = 8'h29;
    mem[12'h4c4] = 8'h33;
    mem[12'h4c5] = 8'h27;
    mem[12'h4c6] = 8'h0a;
    mem[12'h4c7] = 8'h18;
    mem[12'h4c8] = 8'h67;
    mem[12'h4c9] = 8'h29;
    mem[12'h4ca] = 8'h31;
    mem[12'h4cb] = 8'h27;
    mem[12'h4cc] = 8'h0a;
    mem[12'h4cd] = 8'h17;
    mem[12'h4ce] = 8'h69;
    mem[12'h4cf] = 8'h2b;
    mem[12'h4d0] = 8'h2e;
    mem[12'h4d1] = 8'h27;
    mem[12'h4d2] = 8'h0a;
    mem[12'h4d3] = 8'h15;
    mem[12'h4d4] = 8'h6c;
    mem[12'h4d5] = 8'h2d;
    mem[12'h4d6] = 8'h2b;
    mem[12'h4d7] = 8'h27;
    mem[12'h4d8] = 8'h0a;
    mem[12'h4d9] = 8'h14;
    mem[12'h4da] = 8'h6e;
    mem[12'h4db] = 8'h2f;
    mem[12'h4dc] = 8'h28;
    mem[12'h4dd] = 8'h27;
    mem[12'h4de] = 8'h0a;
    mem[12'h4df] = 8'h13;
    mem[12'h4e0] = 8'h71;
    mem[12'h4e1] = 8'h30;
    mem[12'h4e2] = 8'h25;
    mem[12'h4e3] = 8'h27;
    mem[12'h4e4] = 8'h0a;
    mem[12'h4e5] = 8'h11;
    mem[12'h4e6] = 8'h74;
    mem[12'h4e7] = 8'h33;
    mem[12'h4e8] = 8'h21;
    mem[12'h4e9] = 8'h27;
    mem[12'h4ea] = 8'h0a;
    mem[12'h4eb] = 8'h10;
    mem[12'h4ec] = 8'h77;
    mem[12'h4ed] = 8'h36;
    mem[12'h4ee] = 8'h1c;
    mem[12'h4ef] = 8'h27;
    mem[12'h4f0] = 8'h0a;
    mem[12'h4f1] = 8'h0f;
    mem[12'h4f2] = 8'h79;
    mem[12'h4f3] = 8'h3c;
    mem[12'h4f4] = 8'h15;
    mem[12'h4f5] = 8'h27;
    mem[12'h4f6] = 8'h0a;
    mem[12'h4f7] = 8'h0d;
    mem[12'h4f8] = 8'h7d;
    mem[12'h4f9] = 8'h78;
    mem[12'h4fa] = 8'h0a;
    mem[12'h4fb] = 8'h0c;
    mem[12'h4fc] = 8'h7f;
    mem[12'h4fd] = 8'h77;
    mem[12'h4fe] = 8'h0a;
    mem[12'h4ff] = 8'h0a;
    mem[12'h500] = 8'h83;
    mem[12'h501] = 8'h75;
    mem[12'h502] = 8'h0a;
    mem[12'h503] = 8'h08;
    mem[12'h504] = 8'h87;
    mem[12'h505] = 8'h73;
    mem[12'h506] = 8'h0a;
    mem[12'h507] = 8'h07;
    mem[12'h508] = 8'h89;
    mem[12'h509] = 8'h72;
    mem[12'h50a] = 8'h0a;
    mem[12'h50b] = 8'h05;
    mem[12'h50c] = 8'h8d;
    mem[12'h50d] = 8'h70;
    mem[12'h50e] = 8'h0a;
    mem[12'h50f] = 8'h03;
    mem[12'h510] = 8'h91;
    mem[12'h511] = 8'h6e;
    mem[12'h512] = 8'h0a;
    mem[12'h513] = 8'h01;
    mem[12'h514] = 8'h95;
    mem[12'h515] = 8'h6c;
    mem[12'h516] = 8'ha4;
    mem[12'h517] = 8'h6a;
    mem[12'h518] = 8'ha6;
    mem[12'h519] = 8'h68;
    mem[12'h51a] = 8'ha8;
    mem[12'h51b] = 8'h66;
    mem[12'h51c] = 8'hab;
    mem[12'h51d] = 8'h63;
    mem[12'h51e] = 8'had;
    mem[12'h51f] = 8'h61;
    mem[12'h520] = 8'hb0;
    mem[12'h521] = 8'h5b;
    mem[12'h522] = 8'hb6;
    mem[12'h523] = 8'h55;
    mem[12'h524] = 8'hbc;
    mem[12'h525] = 8'h4f;
    mem[12'h526] = 8'hc2;
    mem[12'h527] = 8'h49;
    mem[12'h528] = 8'hc9;
    mem[12'h529] = 8'h41;
    mem[12'h52a] = 8'hd1;
    mem[12'h52b] = 8'h39;
    mem[12'h52c] = 8'hda;
    mem[12'h52d] = 8'h2f;
    mem[12'h52e] = 8'he5;
    mem[12'h52f] = 8'h22;
    mem[12'h530] = 8'hf9;
    mem[12'h531] = 8'h0a;
  end
  assign len = mem[addr];
endmodule
